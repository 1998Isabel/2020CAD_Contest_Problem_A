//
// Conformal-LEC Version 19.20-d218 (25-Feb-2020)
//
module top( C, D, O);
input C, D;
output O;


_DC \n6_5[1] ( O, C, D);

endmodule


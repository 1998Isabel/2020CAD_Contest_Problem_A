//
// Conformal-LEC Version 19.20-d218 (25-Feb-2020)
//
module top(\A[2][9] ,\A[2][8] ,\A[2][7] ,\A[2][6] ,\A[2][5] ,\A[2][4] ,\A[2][3] ,\A[2][2] ,\A[2][1] ,
        \A[2][0] ,\A[1][9] ,\A[1][8] ,\A[1][7] ,\A[1][6] ,\A[1][5] ,\A[1][4] ,\A[1][3] ,\A[1][2] ,\A[1][1] ,
        \A[1][0] ,\A[0][9] ,\A[0][8] ,\A[0][7] ,\A[0][6] ,\A[0][5] ,\A[0][4] ,\A[0][3] ,\A[0][2] ,\A[0][1] ,
        \A[0][0] ,\B[9] ,\B[8] ,\B[7] ,\B[6] ,\B[5] ,\B[4] ,\B[3] ,\B[2] ,\B[1] ,
        \B[0] ,\I[7] ,\I[6] ,\I[5] ,\I[4] ,\I[3] ,\I[2] ,\I[1] ,\I[0] ,\O[19] ,
        \O[18] ,\O[17] ,\O[16] ,\O[15] ,\O[14] ,\O[13] ,\O[12] ,\O[11] ,\O[10] ,\O[9] ,
        \O[8] ,\O[7] ,\O[6] ,\O[5] ,\O[4] ,\O[3] ,\O[2] ,\O[1] ,\O[0] );
input [1:0] \A[2][9] ,\A[2][8] ,\A[2][7] ,\A[2][6] ,\A[2][5] ,\A[2][4] ,\A[2][3] ,\A[2][2] ,\A[2][1] ,        \A[2][0] ,\A[1][9] ,\A[1][8] ,\A[1][7] ,\A[1][6] ,\A[1][5] ,\A[1][4] ,\A[1][3] ,\A[1][2] ,\A[1][1] ,        \A[1][0] ,\A[0][9] ,\A[0][8] ,\A[0][7] ,\A[0][6] ,\A[0][5] ,\A[0][4] ,\A[0][3] ,\A[0][2] ,\A[0][1] ,        \A[0][0] ,\B[9] ,\B[8] ,\B[7] ,\B[6] ,\B[5] ,\B[4] ,\B[3] ,\B[2] ,\B[1] ,        \B[0] ,\I[7] ,\I[6] ,\I[5] ,\I[4] ,\I[3] ,\I[2] ,\I[1] ,\I[0] ;
output [1:0] \O[19] ,\O[18] ,\O[17] ,\O[16] ,\O[15] ,\O[14] ,\O[13] ,\O[12] ,\O[11] ,        \O[10] ,\O[9] ,\O[8] ,\O[7] ,\O[6] ,\O[5] ,\O[4] ,\O[3] ,\O[2] ,\O[1] ,        \O[0] ;

wire [1:0] \69_ZERO , \70_ZERO , \71_ZERO , \72_ZERO , \73_ZERO , \74_ZERO , \75_ZERO , \76 , \77 ,         \78 , \79 , \80 , \81 , \82 , \83 , \84 , \85 , \86_ONE , \87_ONE ,         \88 , \89 , \90 , \91 , \92 , \93 , \94 , \95 , \96 , \97 ,         \98 , \99 , \100 , \101 , \102 , \103 , \104 , \105 , \106 , \107 ,         \108 , \109_A[9] , \110 , \111 , \112 , \113 , \114 , \115_A[8] , \116 , \117 ,         \118 , \119 , \120 , \121_A[7] , \122 , \123 , \124 , \125 , \126 , \127_A[6] ,         \128 , \129 , \130 , \131 , \132 , \133_A[5] , \134 , \135 , \136 , \137 ,         \138 , \139_A[4] , \140 , \141 , \142 , \143 , \144 , \145_A[3] , \146 , \147 ,         \148 , \149 , \150 , \151_A[2] , \152 , \153 , \154 , \155 , \156 , \157_A[1] ,         \158 , \159 , \160 , \161 , \162 , \163_A[0] , \164_B[9] , \165_B[8] , \166_B[7] , \167_B[6] ,         \168_B[5] , \169_B[4] , \170_B[3] , \171_B[2] , \172_B[1] , \173_B[0] , \174 , \175 , \176 , \177 ,         \178 , \179 , \180 , \181 , \182 , \183 , \184 , \185 , \186 , \187 ,         \188 , \189 , \190 , \191 , \192 , \193 , \194 , \195 , \196 , \197 ,         \198 , \199 , \200 , \201 , \202 , \203 , \204 , \205 , \206 , \207 ,         \208 , \209 , \210 , \211 , \212 , \213 , \214 , \215 , \216 , \217 ,         \218 , \219 , \220 , \221 , \222 , \223 , \224 , \225 , \226 , \227 ,         \228 , \229 , \230 , \231 , \232 , \233 , \234 , \235 , \236 , \237 ,         \238 , \239 , \240 , \241 , \242 , \243 , \244 , \245 , \246 , \247 ,         \248 , \249 , \250 , \251 , \252 , \253 , \254 , \255 , \256 , \257 ,         \258 , \259 , \260 , \261 , \262 , \263 , \264 , \265 , \266 , \267 ,         \268 , \269 , \270 , \271 , \272 , \273 , \274 , \275 , \276 , \277 ,         \278 , \279 , \280 , \281 , \282 , \283 , \284 , \285 , \286 , \287 ,         \288 , \289 , \290 , \291 , \292 , \293 , \294 , \295 , \296 , \297 ,         \298 , \299 , \300 , \301 , \302 , \303 , \304 , \305 , \306 , \307 ,         \308 , \309 , \310 , \311 , \312 , \313 , \314 , \315 , \316 , \317 ,         \318 , \319 , \320 , \321 , \322 , \323 , \324 , \325 , \326 , \327 ,         \328 , \329 , \330 , \331 , \332 , \333 , \334 , \335 , \336 , \337 ,         \338 , \339 , \340 , \341 , \342 , \343 , \344 , \345 , \346 , \347 ,         \348 , \349 , \350 , \351 , \352 , \353 , \354 , \355 , \356 , \357 ,         \358 , \359 , \360 , \361 , \362 , \363 , \364 , \365 , \366 , \367 ,         \368 , \369 , \370 , \371 , \372 , \373 , \374 , \375 , \376 , \377 ,         \378 , \379 , \380 , \381 , \382 , \383 , \384 , \385 , \386 , \387 ,         \388 , \389 , \390 , \391 , \392 , \393 , \394 , \395 , \396 , \397 ,         \398 , \399 , \400 , \401 , \402 , \403 , \404 , \405 , \406 , \407 ,         \408 , \409 , \410 , \411 , \412 , \413 , \414 , \415 , \416 , \417 ,         \418 , \419 , \420 , \421 , \422 , \423 , \424 , \425 , \426 , \427 ,         \428 , \429 , \430 , \431 , \432 , \433 , \434 , \435 , \436 , \437 ,         \438 , \439 , \440 , \441 , \442 , \443 , \444 , \445 , \446 , \447 ,         \448 , \449 , \450 , \451 , \452 , \453 , \454 , \455 , \456 , \457 ,         \458 , \459 , \460 , \461 , \462 , \463 , \464 , \465 , \466 , \467 ,         \468 , \469 , \470 , \471 , \472 , \473 , \474 , \475 , \476 , \477 ,         \478 , \479 , \480 , \481 , \482 , \483 , \484 , \485 , \486 , \487 ,         \488 , \489 , \490 , \491 , \492 , \493 , \494 , \495 , \496 , \497 ,         \498 , \499 , \500 , \501 , \502 , \503 , \504 , \505 , \506 , \507 ,         \508 , \509 , \510 , \511 , \512 , \513 , \514 , \515 , \516 , \517 ,         \518 , \519 , \520 , \521 , \522 , \523 , \524 , \525 , \526 , \527 ,         \528 , \529 , \530 , \531 , \532 , \533 , \534 , \535 , \536 , \537 ,         \538 , \539 , \540 , \541 , \542 , \543 , \544 , \545 , \546 , \547 ,         \548 , \549 , \550 , \551 , \552 , \553 , \554 , \555 , \556 , \557 ,         \558 , \559 , \560 , \561 , \562 , \563 , \564 , \565 , \566 , \567 ,         \568 , \569 , \570 , \571 , \572 , \573 , \574 , \575 , \576 , \577 ,         \578 , \579 , \580 , \581 , \582 , \583 , \584 , \585 , \586 , \587 ,         \588 , \589 , \590 , \591 , \592 , \593 , \594 , \595 , \596 , \597 ,         \598 , \599 , \600 , \601 , \602 , \603 , \604 , \605 , \606 , \607 ,         \608 , \609 , \610 , \611 , \612 , \613 , \614 , \615 , \616 , \617 ,         \618 , \619 , \620 , \621 , \622 , \623 , \624 , \625 , \626 , \627 ,         \628 , \629 , \630 , \631 , \632 , \633 , \634 , \635 , \636 , \637 ,         \638 , \639 , \640 , \641 , \642 , \643 , \644 , \645 , \646 , \647 ,         \648 , \649 , \650 , \651 , \652 , \653 , \654 , \655 , \656 , \657 ,         \658 , \659 , \660 , \661 , \662 , \663 , \664 , \665 , \666 , \667 ,         \668 , \669 , \670 , \671 , \672 , \673 , \674 , \675_Z[19] , \676 , \677_Z[18] ,         \678 , \679_Z[17] , \680 , \681_Z[16] , \682 , \683_Z[15] , \684 , \685_Z[14] , \686 , \687_Z[13] ,         \688 , \689_Z[12] , \690 , \691_Z[11] , \692 , \693_Z[10] , \694 , \695_Z[9] , \696 , \697_Z[8] ,         \698 , \699_Z[7] , \700 , \701_Z[6] , \702 , \703_Z[5] , \704 , \705_Z[4] , \706 , \707_Z[3] ,         \708 , \709_Z[2] , \710 , \711_Z[1] , \712 , \713_Z[0] ;
mbuf \U$labaj85 ( \O[19] , \675_Z[19] );
mbuf \U$labaj86 ( \O[18] , \677_Z[18] );
mbuf \U$labaj87 ( \O[17] , \679_Z[17] );
mbuf \U$labaj88 ( \O[16] , \681_Z[16] );
mbuf \U$labaj89 ( \O[15] , \683_Z[15] );
mbuf \U$labaj90 ( \O[14] , \685_Z[14] );
mbuf \U$labaj91 ( \O[13] , \687_Z[13] );
mbuf \U$labaj92 ( \O[12] , \689_Z[12] );
mbuf \U$labaj93 ( \O[11] , \691_Z[11] );
mbuf \U$labaj94 ( \O[10] , \693_Z[10] );
mbuf \U$labaj95 ( \O[9] , \695_Z[9] );
mbuf \U$labaj96 ( \O[8] , \697_Z[8] );
mbuf \U$labaj97 ( \O[7] , \699_Z[7] );
mbuf \U$labaj98 ( \O[6] , \701_Z[6] );
mbuf \U$labaj99 ( \O[5] , \703_Z[5] );
mbuf \U$labaj100 ( \O[4] , \705_Z[4] );
mbuf \U$labaj101 ( \O[3] , \707_Z[3] );
mbuf \U$labaj102 ( \O[2] , \709_Z[2] );
mbuf \U$labaj103 ( \O[1] , \711_Z[1] );
mbuf \U$labaj104 ( \O[0] , \713_Z[0] );
mnot \U$7 ( \88 , \I[1] );
mnor \U$8 ( \89 , \I[0] , \88 , \I[2] , \I[3] , \I[4] , \I[5] , \I[6] , \I[7] );
mand \U$3/U$40 ( \90 , \A[2][9] , \89 );
mnot \U$5 ( \91 , \I[0] );
mnor \U$6 ( \92 , \91 , \I[1] , \I[2] , \I[3] , \I[4] , \I[5] , \I[6] , \I[7] );
mand \U$3/U$39 ( \93 , \A[1][9] , \92 );
mnor \U$4 ( \94 , \I[0] , \I[1] , \I[2] , \I[3] , \I[4] , \I[5] , \I[6] , \I[7] );
mand \U$3/U$38 ( \95 , \A[0][9] , \94 );
mor \U$3/U$37 ( \96 , \90 , \93 , \95 );
mbuf \U$2/A[2] ( \97 , \I[2] );
mbuf \U$2/A[3] ( \98 , \I[3] );
mbuf \U$2/A[4] ( \99 , \I[4] );
mbuf \U$2/A[5] ( \100 , \I[5] );
mbuf \U$2/A[6] ( \101 , \I[6] );
mbuf \U$2/A[7] ( \102 , \I[7] );
mbuf \U$2/A[1] ( \103 , \I[1] );
mbuf \U$2/A[0] ( \104 , \I[0] );
mand \U$2/U$2 ( \105 , \103 , \104 );
mor \U$2/U$1 ( \106 , \97 , \98 , \99 , \100 , \101 , \102 , \105 );
mbuf \U$2/Z ( \107 , \106 );
m_DC \n6_5[9] ( \108 , \96 , \107 );
mbuf \mul_6_19/A[9] ( \109_A[9] , \108 );
mand \U$3/U$36 ( \110 , \A[2][8] , \89 );
mand \U$3/U$35 ( \111 , \A[1][8] , \92 );
mand \U$3/U$34 ( \112 , \A[0][8] , \94 );
mor \U$3/U$33 ( \113 , \110 , \111 , \112 );
m_DC \n6_5[8] ( \114 , \113 , \107 );
mbuf \mul_6_19/A[8] ( \115_A[8] , \114 );
mand \U$3/U$32 ( \116 , \A[2][7] , \89 );
mand \U$3/U$31 ( \117 , \A[1][7] , \92 );
mand \U$3/U$30 ( \118 , \A[0][7] , \94 );
mor \U$3/U$29 ( \119 , \116 , \117 , \118 );
m_DC \n6_5[7] ( \120 , \119 , \107 );
mbuf \mul_6_19/A[7] ( \121_A[7] , \120 );
mand \U$3/U$28 ( \122 , \A[2][6] , \89 );
mand \U$3/U$27 ( \123 , \A[1][6] , \92 );
mand \U$3/U$26 ( \124 , \A[0][6] , \94 );
mor \U$3/U$25 ( \125 , \122 , \123 , \124 );
m_DC \n6_5[6] ( \126 , \125 , \107 );
mbuf \mul_6_19/A[6] ( \127_A[6] , \126 );
mand \U$3/U$24 ( \128 , \A[2][5] , \89 );
mand \U$3/U$23 ( \129 , \A[1][5] , \92 );
mand \U$3/U$22 ( \130 , \A[0][5] , \94 );
mor \U$3/U$21 ( \131 , \128 , \129 , \130 );
m_DC \n6_5[5] ( \132 , \131 , \107 );
mbuf \mul_6_19/A[5] ( \133_A[5] , \132 );
mand \U$3/U$20 ( \134 , \A[2][4] , \89 );
mand \U$3/U$19 ( \135 , \A[1][4] , \92 );
mand \U$3/U$18 ( \136 , \A[0][4] , \94 );
mor \U$3/U$17 ( \137 , \134 , \135 , \136 );
m_DC \n6_5[4] ( \138 , \137 , \107 );
mbuf \mul_6_19/A[4] ( \139_A[4] , \138 );
mand \U$3/U$16 ( \140 , \A[2][3] , \89 );
mand \U$3/U$15 ( \141 , \A[1][3] , \92 );
mand \U$3/U$14 ( \142 , \A[0][3] , \94 );
mor \U$3/U$13 ( \143 , \140 , \141 , \142 );
m_DC \n6_5[3] ( \144 , \143 , \107 );
mbuf \mul_6_19/A[3] ( \145_A[3] , \144 );
mand \U$3/U$12 ( \146 , \A[2][2] , \89 );
mand \U$3/U$11 ( \147 , \A[1][2] , \92 );
mand \U$3/U$10 ( \148 , \A[0][2] , \94 );
mor \U$3/U$9 ( \149 , \146 , \147 , \148 );
m_DC \n6_5[2] ( \150 , \149 , \107 );
mbuf \mul_6_19/A[2] ( \151_A[2] , \150 );
mand \U$3/U$8 ( \152 , \A[2][1] , \89 );
mand \U$3/U$7 ( \153 , \A[1][1] , \92 );
mand \U$3/U$6 ( \154 , \A[0][1] , \94 );
mor \U$3/U$5 ( \155 , \152 , \153 , \154 );
m_DC \n6_5[1] ( \156 , \155 , \107 );
mbuf \mul_6_19/A[1] ( \157_A[1] , \156 );
mand \U$3/U$4 ( \158 , \A[2][0] , \89 );
mand \U$3/U$3 ( \159 , \A[1][0] , \92 );
mand \U$3/U$2 ( \160 , \A[0][0] , \94 );
mor \U$3/U$1 ( \161 , \158 , \159 , \160 );
m_DC \n6_5[0] ( \162 , \161 , \107 );
mbuf \mul_6_19/A[0] ( \163_A[0] , \162 );
mbuf \mul_6_19/B[9] ( \164_B[9] , \B[9] );
mbuf \mul_6_19/B[8] ( \165_B[8] , \B[8] );
mbuf \mul_6_19/B[7] ( \166_B[7] , \B[7] );
mbuf \mul_6_19/B[6] ( \167_B[6] , \B[6] );
mbuf \mul_6_19/B[5] ( \168_B[5] , \B[5] );
mbuf \mul_6_19/B[4] ( \169_B[4] , \B[4] );
mbuf \mul_6_19/B[3] ( \170_B[3] , \B[3] );
mbuf \mul_6_19/B[2] ( \171_B[2] , \B[2] );
mbuf \mul_6_19/B[1] ( \172_B[1] , \B[1] );
mbuf \mul_6_19/B[0] ( \173_B[0] , \B[0] );
mand \mul_6_19/U$501 ( \174 , \109_A[9] , \172_B[1] );
mand \mul_6_19/U$511 ( \175 , \109_A[9] , \173_B[0] );
mand \mul_6_19/U$502 ( \176 , \115_A[8] , \172_B[1] );
mand \mul_6_19/U$462 ( \177 , \175 , \176 );
mxor \mul_6_19/U$463 ( \178 , \175 , \176 );
mand \mul_6_19/U$512 ( \179 , \115_A[8] , \173_B[0] );
mand \mul_6_19/U$503 ( \180 , \121_A[7] , \172_B[1] );
mand \mul_6_19/U$467 ( \181 , \179 , \180 );
mxor \mul_6_19/U$468 ( \182 , \179 , \180 );
mand \mul_6_19/U$513 ( \183 , \121_A[7] , \173_B[0] );
mand \mul_6_19/U$504 ( \184 , \127_A[6] , \172_B[1] );
mand \mul_6_19/U$472 ( \185 , \183 , \184 );
mxor \mul_6_19/U$473 ( \186 , \183 , \184 );
mand \mul_6_19/U$514 ( \187 , \127_A[6] , \173_B[0] );
mand \mul_6_19/U$505 ( \188 , \133_A[5] , \172_B[1] );
mand \mul_6_19/U$477 ( \189 , \187 , \188 );
mxor \mul_6_19/U$478 ( \190 , \187 , \188 );
mand \mul_6_19/U$515 ( \191 , \133_A[5] , \173_B[0] );
mand \mul_6_19/U$506 ( \192 , \139_A[4] , \172_B[1] );
mand \mul_6_19/U$482 ( \193 , \191 , \192 );
mxor \mul_6_19/U$483 ( \194 , \191 , \192 );
mand \mul_6_19/U$516 ( \195 , \139_A[4] , \173_B[0] );
mand \mul_6_19/U$507 ( \196 , \145_A[3] , \172_B[1] );
mand \mul_6_19/U$487 ( \197 , \195 , \196 );
mxor \mul_6_19/U$488 ( \198 , \195 , \196 );
mand \mul_6_19/U$517 ( \199 , \145_A[3] , \173_B[0] );
mand \mul_6_19/U$508 ( \200 , \151_A[2] , \172_B[1] );
mand \mul_6_19/U$492 ( \201 , \199 , \200 );
mxor \mul_6_19/U$493 ( \202 , \199 , \200 );
mand \mul_6_19/U$518 ( \203 , \151_A[2] , \173_B[0] );
mand \mul_6_19/U$509 ( \204 , \157_A[1] , \172_B[1] );
mand \mul_6_19/U$497 ( \205 , \203 , \204 );
mxor \mul_6_19/U$498 ( \206 , \203 , \204 );
mand \mul_6_19/U$519 ( \207 , \157_A[1] , \173_B[0] );
mand \mul_6_19/U$510 ( \208 , \163_A[0] , \172_B[1] );
mand \mul_6_19/U$499 ( \209 , \207 , \208 );
mand \mul_6_19/U$496 ( \210 , \206 , \209 );
mor \mul_6_19/U$494 ( \211 , \205 , \210 );
mand \mul_6_19/U$491 ( \212 , \202 , \211 );
mor \mul_6_19/U$489 ( \213 , \201 , \212 );
mand \mul_6_19/U$486 ( \214 , \198 , \213 );
mor \mul_6_19/U$484 ( \215 , \197 , \214 );
mand \mul_6_19/U$481 ( \216 , \194 , \215 );
mor \mul_6_19/U$479 ( \217 , \193 , \216 );
mand \mul_6_19/U$476 ( \218 , \190 , \217 );
mor \mul_6_19/U$474 ( \219 , \189 , \218 );
mand \mul_6_19/U$471 ( \220 , \186 , \219 );
mor \mul_6_19/U$469 ( \221 , \185 , \220 );
mand \mul_6_19/U$466 ( \222 , \182 , \221 );
mor \mul_6_19/U$464 ( \223 , \181 , \222 );
mand \mul_6_19/U$461 ( \224 , \178 , \223 );
mor \mul_6_19/U$459 ( \225 , \177 , \224 );
mand \mul_6_19/U$458 ( \226 , \174 , \225 );
mand \mul_6_19/U$447 ( \227 , \109_A[9] , \171_B[2] );
mand \mul_6_19/U$403 ( \228 , \226 , \227 );
mxor \mul_6_19/U$404 ( \229 , \226 , \227 );
mxor \mul_6_19/U$457 ( \230 , \174 , \225 );
mand \mul_6_19/U$448 ( \231 , \115_A[8] , \171_B[2] );
mand \mul_6_19/U$408 ( \232 , \230 , \231 );
mxor \mul_6_19/U$409 ( \233 , \230 , \231 );
mxor \mul_6_19/U$460 ( \234 , \178 , \223 );
mand \mul_6_19/U$449 ( \235 , \121_A[7] , \171_B[2] );
mand \mul_6_19/U$413 ( \236 , \234 , \235 );
mxor \mul_6_19/U$414 ( \237 , \234 , \235 );
mxor \mul_6_19/U$465 ( \238 , \182 , \221 );
mand \mul_6_19/U$450 ( \239 , \127_A[6] , \171_B[2] );
mand \mul_6_19/U$418 ( \240 , \238 , \239 );
mxor \mul_6_19/U$419 ( \241 , \238 , \239 );
mxor \mul_6_19/U$470 ( \242 , \186 , \219 );
mand \mul_6_19/U$451 ( \243 , \133_A[5] , \171_B[2] );
mand \mul_6_19/U$423 ( \244 , \242 , \243 );
mxor \mul_6_19/U$424 ( \245 , \242 , \243 );
mxor \mul_6_19/U$475 ( \246 , \190 , \217 );
mand \mul_6_19/U$452 ( \247 , \139_A[4] , \171_B[2] );
mand \mul_6_19/U$428 ( \248 , \246 , \247 );
mxor \mul_6_19/U$429 ( \249 , \246 , \247 );
mxor \mul_6_19/U$480 ( \250 , \194 , \215 );
mand \mul_6_19/U$453 ( \251 , \145_A[3] , \171_B[2] );
mand \mul_6_19/U$433 ( \252 , \250 , \251 );
mxor \mul_6_19/U$434 ( \253 , \250 , \251 );
mxor \mul_6_19/U$485 ( \254 , \198 , \213 );
mand \mul_6_19/U$454 ( \255 , \151_A[2] , \171_B[2] );
mand \mul_6_19/U$438 ( \256 , \254 , \255 );
mxor \mul_6_19/U$439 ( \257 , \254 , \255 );
mxor \mul_6_19/U$490 ( \258 , \202 , \211 );
mand \mul_6_19/U$455 ( \259 , \157_A[1] , \171_B[2] );
mand \mul_6_19/U$443 ( \260 , \258 , \259 );
mxor \mul_6_19/U$444 ( \261 , \258 , \259 );
mxor \mul_6_19/U$495 ( \262 , \206 , \209 );
mand \mul_6_19/U$456 ( \263 , \163_A[0] , \171_B[2] );
mand \mul_6_19/U$445 ( \264 , \262 , \263 );
mand \mul_6_19/U$442 ( \265 , \261 , \264 );
mor \mul_6_19/U$440 ( \266 , \260 , \265 );
mand \mul_6_19/U$437 ( \267 , \257 , \266 );
mor \mul_6_19/U$435 ( \268 , \256 , \267 );
mand \mul_6_19/U$432 ( \269 , \253 , \268 );
mor \mul_6_19/U$430 ( \270 , \252 , \269 );
mand \mul_6_19/U$427 ( \271 , \249 , \270 );
mor \mul_6_19/U$425 ( \272 , \248 , \271 );
mand \mul_6_19/U$422 ( \273 , \245 , \272 );
mor \mul_6_19/U$420 ( \274 , \244 , \273 );
mand \mul_6_19/U$417 ( \275 , \241 , \274 );
mor \mul_6_19/U$415 ( \276 , \240 , \275 );
mand \mul_6_19/U$412 ( \277 , \237 , \276 );
mor \mul_6_19/U$410 ( \278 , \236 , \277 );
mand \mul_6_19/U$407 ( \279 , \233 , \278 );
mor \mul_6_19/U$405 ( \280 , \232 , \279 );
mand \mul_6_19/U$402 ( \281 , \229 , \280 );
mor \mul_6_19/U$400 ( \282 , \228 , \281 );
mand \mul_6_19/U$390 ( \283 , \109_A[9] , \170_B[3] );
mand \mul_6_19/U$346 ( \284 , \282 , \283 );
mxor \mul_6_19/U$347 ( \285 , \282 , \283 );
mxor \mul_6_19/U$401 ( \286 , \229 , \280 );
mand \mul_6_19/U$391 ( \287 , \115_A[8] , \170_B[3] );
mand \mul_6_19/U$351 ( \288 , \286 , \287 );
mxor \mul_6_19/U$352 ( \289 , \286 , \287 );
mxor \mul_6_19/U$406 ( \290 , \233 , \278 );
mand \mul_6_19/U$392 ( \291 , \121_A[7] , \170_B[3] );
mand \mul_6_19/U$356 ( \292 , \290 , \291 );
mxor \mul_6_19/U$357 ( \293 , \290 , \291 );
mxor \mul_6_19/U$411 ( \294 , \237 , \276 );
mand \mul_6_19/U$393 ( \295 , \127_A[6] , \170_B[3] );
mand \mul_6_19/U$361 ( \296 , \294 , \295 );
mxor \mul_6_19/U$362 ( \297 , \294 , \295 );
mxor \mul_6_19/U$416 ( \298 , \241 , \274 );
mand \mul_6_19/U$394 ( \299 , \133_A[5] , \170_B[3] );
mand \mul_6_19/U$366 ( \300 , \298 , \299 );
mxor \mul_6_19/U$367 ( \301 , \298 , \299 );
mxor \mul_6_19/U$421 ( \302 , \245 , \272 );
mand \mul_6_19/U$395 ( \303 , \139_A[4] , \170_B[3] );
mand \mul_6_19/U$371 ( \304 , \302 , \303 );
mxor \mul_6_19/U$372 ( \305 , \302 , \303 );
mxor \mul_6_19/U$426 ( \306 , \249 , \270 );
mand \mul_6_19/U$396 ( \307 , \145_A[3] , \170_B[3] );
mand \mul_6_19/U$376 ( \308 , \306 , \307 );
mxor \mul_6_19/U$377 ( \309 , \306 , \307 );
mxor \mul_6_19/U$431 ( \310 , \253 , \268 );
mand \mul_6_19/U$397 ( \311 , \151_A[2] , \170_B[3] );
mand \mul_6_19/U$381 ( \312 , \310 , \311 );
mxor \mul_6_19/U$382 ( \313 , \310 , \311 );
mxor \mul_6_19/U$436 ( \314 , \257 , \266 );
mand \mul_6_19/U$398 ( \315 , \157_A[1] , \170_B[3] );
mand \mul_6_19/U$386 ( \316 , \314 , \315 );
mxor \mul_6_19/U$387 ( \317 , \314 , \315 );
mxor \mul_6_19/U$441 ( \318 , \261 , \264 );
mand \mul_6_19/U$399 ( \319 , \163_A[0] , \170_B[3] );
mand \mul_6_19/U$388 ( \320 , \318 , \319 );
mand \mul_6_19/U$385 ( \321 , \317 , \320 );
mor \mul_6_19/U$383 ( \322 , \316 , \321 );
mand \mul_6_19/U$380 ( \323 , \313 , \322 );
mor \mul_6_19/U$378 ( \324 , \312 , \323 );
mand \mul_6_19/U$375 ( \325 , \309 , \324 );
mor \mul_6_19/U$373 ( \326 , \308 , \325 );
mand \mul_6_19/U$370 ( \327 , \305 , \326 );
mor \mul_6_19/U$368 ( \328 , \304 , \327 );
mand \mul_6_19/U$365 ( \329 , \301 , \328 );
mor \mul_6_19/U$363 ( \330 , \300 , \329 );
mand \mul_6_19/U$360 ( \331 , \297 , \330 );
mor \mul_6_19/U$358 ( \332 , \296 , \331 );
mand \mul_6_19/U$355 ( \333 , \293 , \332 );
mor \mul_6_19/U$353 ( \334 , \292 , \333 );
mand \mul_6_19/U$350 ( \335 , \289 , \334 );
mor \mul_6_19/U$348 ( \336 , \288 , \335 );
mand \mul_6_19/U$345 ( \337 , \285 , \336 );
mor \mul_6_19/U$343 ( \338 , \284 , \337 );
mand \mul_6_19/U$333 ( \339 , \109_A[9] , \169_B[4] );
mand \mul_6_19/U$289 ( \340 , \338 , \339 );
mxor \mul_6_19/U$290 ( \341 , \338 , \339 );
mxor \mul_6_19/U$344 ( \342 , \285 , \336 );
mand \mul_6_19/U$334 ( \343 , \115_A[8] , \169_B[4] );
mand \mul_6_19/U$294 ( \344 , \342 , \343 );
mxor \mul_6_19/U$295 ( \345 , \342 , \343 );
mxor \mul_6_19/U$349 ( \346 , \289 , \334 );
mand \mul_6_19/U$335 ( \347 , \121_A[7] , \169_B[4] );
mand \mul_6_19/U$299 ( \348 , \346 , \347 );
mxor \mul_6_19/U$300 ( \349 , \346 , \347 );
mxor \mul_6_19/U$354 ( \350 , \293 , \332 );
mand \mul_6_19/U$336 ( \351 , \127_A[6] , \169_B[4] );
mand \mul_6_19/U$304 ( \352 , \350 , \351 );
mxor \mul_6_19/U$305 ( \353 , \350 , \351 );
mxor \mul_6_19/U$359 ( \354 , \297 , \330 );
mand \mul_6_19/U$337 ( \355 , \133_A[5] , \169_B[4] );
mand \mul_6_19/U$309 ( \356 , \354 , \355 );
mxor \mul_6_19/U$310 ( \357 , \354 , \355 );
mxor \mul_6_19/U$364 ( \358 , \301 , \328 );
mand \mul_6_19/U$338 ( \359 , \139_A[4] , \169_B[4] );
mand \mul_6_19/U$314 ( \360 , \358 , \359 );
mxor \mul_6_19/U$315 ( \361 , \358 , \359 );
mxor \mul_6_19/U$369 ( \362 , \305 , \326 );
mand \mul_6_19/U$339 ( \363 , \145_A[3] , \169_B[4] );
mand \mul_6_19/U$319 ( \364 , \362 , \363 );
mxor \mul_6_19/U$320 ( \365 , \362 , \363 );
mxor \mul_6_19/U$374 ( \366 , \309 , \324 );
mand \mul_6_19/U$340 ( \367 , \151_A[2] , \169_B[4] );
mand \mul_6_19/U$324 ( \368 , \366 , \367 );
mxor \mul_6_19/U$325 ( \369 , \366 , \367 );
mxor \mul_6_19/U$379 ( \370 , \313 , \322 );
mand \mul_6_19/U$341 ( \371 , \157_A[1] , \169_B[4] );
mand \mul_6_19/U$329 ( \372 , \370 , \371 );
mxor \mul_6_19/U$330 ( \373 , \370 , \371 );
mxor \mul_6_19/U$384 ( \374 , \317 , \320 );
mand \mul_6_19/U$342 ( \375 , \163_A[0] , \169_B[4] );
mand \mul_6_19/U$331 ( \376 , \374 , \375 );
mand \mul_6_19/U$328 ( \377 , \373 , \376 );
mor \mul_6_19/U$326 ( \378 , \372 , \377 );
mand \mul_6_19/U$323 ( \379 , \369 , \378 );
mor \mul_6_19/U$321 ( \380 , \368 , \379 );
mand \mul_6_19/U$318 ( \381 , \365 , \380 );
mor \mul_6_19/U$316 ( \382 , \364 , \381 );
mand \mul_6_19/U$313 ( \383 , \361 , \382 );
mor \mul_6_19/U$311 ( \384 , \360 , \383 );
mand \mul_6_19/U$308 ( \385 , \357 , \384 );
mor \mul_6_19/U$306 ( \386 , \356 , \385 );
mand \mul_6_19/U$303 ( \387 , \353 , \386 );
mor \mul_6_19/U$301 ( \388 , \352 , \387 );
mand \mul_6_19/U$298 ( \389 , \349 , \388 );
mor \mul_6_19/U$296 ( \390 , \348 , \389 );
mand \mul_6_19/U$293 ( \391 , \345 , \390 );
mor \mul_6_19/U$291 ( \392 , \344 , \391 );
mand \mul_6_19/U$288 ( \393 , \341 , \392 );
mor \mul_6_19/U$286 ( \394 , \340 , \393 );
mand \mul_6_19/U$276 ( \395 , \109_A[9] , \168_B[5] );
mand \mul_6_19/U$232 ( \396 , \394 , \395 );
mxor \mul_6_19/U$233 ( \397 , \394 , \395 );
mxor \mul_6_19/U$287 ( \398 , \341 , \392 );
mand \mul_6_19/U$277 ( \399 , \115_A[8] , \168_B[5] );
mand \mul_6_19/U$237 ( \400 , \398 , \399 );
mxor \mul_6_19/U$238 ( \401 , \398 , \399 );
mxor \mul_6_19/U$292 ( \402 , \345 , \390 );
mand \mul_6_19/U$278 ( \403 , \121_A[7] , \168_B[5] );
mand \mul_6_19/U$242 ( \404 , \402 , \403 );
mxor \mul_6_19/U$243 ( \405 , \402 , \403 );
mxor \mul_6_19/U$297 ( \406 , \349 , \388 );
mand \mul_6_19/U$279 ( \407 , \127_A[6] , \168_B[5] );
mand \mul_6_19/U$247 ( \408 , \406 , \407 );
mxor \mul_6_19/U$248 ( \409 , \406 , \407 );
mxor \mul_6_19/U$302 ( \410 , \353 , \386 );
mand \mul_6_19/U$280 ( \411 , \133_A[5] , \168_B[5] );
mand \mul_6_19/U$252 ( \412 , \410 , \411 );
mxor \mul_6_19/U$253 ( \413 , \410 , \411 );
mxor \mul_6_19/U$307 ( \414 , \357 , \384 );
mand \mul_6_19/U$281 ( \415 , \139_A[4] , \168_B[5] );
mand \mul_6_19/U$257 ( \416 , \414 , \415 );
mxor \mul_6_19/U$258 ( \417 , \414 , \415 );
mxor \mul_6_19/U$312 ( \418 , \361 , \382 );
mand \mul_6_19/U$282 ( \419 , \145_A[3] , \168_B[5] );
mand \mul_6_19/U$262 ( \420 , \418 , \419 );
mxor \mul_6_19/U$263 ( \421 , \418 , \419 );
mxor \mul_6_19/U$317 ( \422 , \365 , \380 );
mand \mul_6_19/U$283 ( \423 , \151_A[2] , \168_B[5] );
mand \mul_6_19/U$267 ( \424 , \422 , \423 );
mxor \mul_6_19/U$268 ( \425 , \422 , \423 );
mxor \mul_6_19/U$322 ( \426 , \369 , \378 );
mand \mul_6_19/U$284 ( \427 , \157_A[1] , \168_B[5] );
mand \mul_6_19/U$272 ( \428 , \426 , \427 );
mxor \mul_6_19/U$273 ( \429 , \426 , \427 );
mxor \mul_6_19/U$327 ( \430 , \373 , \376 );
mand \mul_6_19/U$285 ( \431 , \163_A[0] , \168_B[5] );
mand \mul_6_19/U$274 ( \432 , \430 , \431 );
mand \mul_6_19/U$271 ( \433 , \429 , \432 );
mor \mul_6_19/U$269 ( \434 , \428 , \433 );
mand \mul_6_19/U$266 ( \435 , \425 , \434 );
mor \mul_6_19/U$264 ( \436 , \424 , \435 );
mand \mul_6_19/U$261 ( \437 , \421 , \436 );
mor \mul_6_19/U$259 ( \438 , \420 , \437 );
mand \mul_6_19/U$256 ( \439 , \417 , \438 );
mor \mul_6_19/U$254 ( \440 , \416 , \439 );
mand \mul_6_19/U$251 ( \441 , \413 , \440 );
mor \mul_6_19/U$249 ( \442 , \412 , \441 );
mand \mul_6_19/U$246 ( \443 , \409 , \442 );
mor \mul_6_19/U$244 ( \444 , \408 , \443 );
mand \mul_6_19/U$241 ( \445 , \405 , \444 );
mor \mul_6_19/U$239 ( \446 , \404 , \445 );
mand \mul_6_19/U$236 ( \447 , \401 , \446 );
mor \mul_6_19/U$234 ( \448 , \400 , \447 );
mand \mul_6_19/U$231 ( \449 , \397 , \448 );
mor \mul_6_19/U$229 ( \450 , \396 , \449 );
mand \mul_6_19/U$219 ( \451 , \109_A[9] , \167_B[6] );
mand \mul_6_19/U$175 ( \452 , \450 , \451 );
mxor \mul_6_19/U$176 ( \453 , \450 , \451 );
mxor \mul_6_19/U$230 ( \454 , \397 , \448 );
mand \mul_6_19/U$220 ( \455 , \115_A[8] , \167_B[6] );
mand \mul_6_19/U$180 ( \456 , \454 , \455 );
mxor \mul_6_19/U$181 ( \457 , \454 , \455 );
mxor \mul_6_19/U$235 ( \458 , \401 , \446 );
mand \mul_6_19/U$221 ( \459 , \121_A[7] , \167_B[6] );
mand \mul_6_19/U$185 ( \460 , \458 , \459 );
mxor \mul_6_19/U$186 ( \461 , \458 , \459 );
mxor \mul_6_19/U$240 ( \462 , \405 , \444 );
mand \mul_6_19/U$222 ( \463 , \127_A[6] , \167_B[6] );
mand \mul_6_19/U$190 ( \464 , \462 , \463 );
mxor \mul_6_19/U$191 ( \465 , \462 , \463 );
mxor \mul_6_19/U$245 ( \466 , \409 , \442 );
mand \mul_6_19/U$223 ( \467 , \133_A[5] , \167_B[6] );
mand \mul_6_19/U$195 ( \468 , \466 , \467 );
mxor \mul_6_19/U$196 ( \469 , \466 , \467 );
mxor \mul_6_19/U$250 ( \470 , \413 , \440 );
mand \mul_6_19/U$224 ( \471 , \139_A[4] , \167_B[6] );
mand \mul_6_19/U$200 ( \472 , \470 , \471 );
mxor \mul_6_19/U$201 ( \473 , \470 , \471 );
mxor \mul_6_19/U$255 ( \474 , \417 , \438 );
mand \mul_6_19/U$225 ( \475 , \145_A[3] , \167_B[6] );
mand \mul_6_19/U$205 ( \476 , \474 , \475 );
mxor \mul_6_19/U$206 ( \477 , \474 , \475 );
mxor \mul_6_19/U$260 ( \478 , \421 , \436 );
mand \mul_6_19/U$226 ( \479 , \151_A[2] , \167_B[6] );
mand \mul_6_19/U$210 ( \480 , \478 , \479 );
mxor \mul_6_19/U$211 ( \481 , \478 , \479 );
mxor \mul_6_19/U$265 ( \482 , \425 , \434 );
mand \mul_6_19/U$227 ( \483 , \157_A[1] , \167_B[6] );
mand \mul_6_19/U$215 ( \484 , \482 , \483 );
mxor \mul_6_19/U$216 ( \485 , \482 , \483 );
mxor \mul_6_19/U$270 ( \486 , \429 , \432 );
mand \mul_6_19/U$228 ( \487 , \163_A[0] , \167_B[6] );
mand \mul_6_19/U$217 ( \488 , \486 , \487 );
mand \mul_6_19/U$214 ( \489 , \485 , \488 );
mor \mul_6_19/U$212 ( \490 , \484 , \489 );
mand \mul_6_19/U$209 ( \491 , \481 , \490 );
mor \mul_6_19/U$207 ( \492 , \480 , \491 );
mand \mul_6_19/U$204 ( \493 , \477 , \492 );
mor \mul_6_19/U$202 ( \494 , \476 , \493 );
mand \mul_6_19/U$199 ( \495 , \473 , \494 );
mor \mul_6_19/U$197 ( \496 , \472 , \495 );
mand \mul_6_19/U$194 ( \497 , \469 , \496 );
mor \mul_6_19/U$192 ( \498 , \468 , \497 );
mand \mul_6_19/U$189 ( \499 , \465 , \498 );
mor \mul_6_19/U$187 ( \500 , \464 , \499 );
mand \mul_6_19/U$184 ( \501 , \461 , \500 );
mor \mul_6_19/U$182 ( \502 , \460 , \501 );
mand \mul_6_19/U$179 ( \503 , \457 , \502 );
mor \mul_6_19/U$177 ( \504 , \456 , \503 );
mand \mul_6_19/U$174 ( \505 , \453 , \504 );
mor \mul_6_19/U$172 ( \506 , \452 , \505 );
mand \mul_6_19/U$162 ( \507 , \109_A[9] , \166_B[7] );
mand \mul_6_19/U$118 ( \508 , \506 , \507 );
mxor \mul_6_19/U$119 ( \509 , \506 , \507 );
mxor \mul_6_19/U$173 ( \510 , \453 , \504 );
mand \mul_6_19/U$163 ( \511 , \115_A[8] , \166_B[7] );
mand \mul_6_19/U$123 ( \512 , \510 , \511 );
mxor \mul_6_19/U$124 ( \513 , \510 , \511 );
mxor \mul_6_19/U$178 ( \514 , \457 , \502 );
mand \mul_6_19/U$164 ( \515 , \121_A[7] , \166_B[7] );
mand \mul_6_19/U$128 ( \516 , \514 , \515 );
mxor \mul_6_19/U$129 ( \517 , \514 , \515 );
mxor \mul_6_19/U$183 ( \518 , \461 , \500 );
mand \mul_6_19/U$165 ( \519 , \127_A[6] , \166_B[7] );
mand \mul_6_19/U$133 ( \520 , \518 , \519 );
mxor \mul_6_19/U$134 ( \521 , \518 , \519 );
mxor \mul_6_19/U$188 ( \522 , \465 , \498 );
mand \mul_6_19/U$166 ( \523 , \133_A[5] , \166_B[7] );
mand \mul_6_19/U$138 ( \524 , \522 , \523 );
mxor \mul_6_19/U$139 ( \525 , \522 , \523 );
mxor \mul_6_19/U$193 ( \526 , \469 , \496 );
mand \mul_6_19/U$167 ( \527 , \139_A[4] , \166_B[7] );
mand \mul_6_19/U$143 ( \528 , \526 , \527 );
mxor \mul_6_19/U$144 ( \529 , \526 , \527 );
mxor \mul_6_19/U$198 ( \530 , \473 , \494 );
mand \mul_6_19/U$168 ( \531 , \145_A[3] , \166_B[7] );
mand \mul_6_19/U$148 ( \532 , \530 , \531 );
mxor \mul_6_19/U$149 ( \533 , \530 , \531 );
mxor \mul_6_19/U$203 ( \534 , \477 , \492 );
mand \mul_6_19/U$169 ( \535 , \151_A[2] , \166_B[7] );
mand \mul_6_19/U$153 ( \536 , \534 , \535 );
mxor \mul_6_19/U$154 ( \537 , \534 , \535 );
mxor \mul_6_19/U$208 ( \538 , \481 , \490 );
mand \mul_6_19/U$170 ( \539 , \157_A[1] , \166_B[7] );
mand \mul_6_19/U$158 ( \540 , \538 , \539 );
mxor \mul_6_19/U$159 ( \541 , \538 , \539 );
mxor \mul_6_19/U$213 ( \542 , \485 , \488 );
mand \mul_6_19/U$171 ( \543 , \163_A[0] , \166_B[7] );
mand \mul_6_19/U$160 ( \544 , \542 , \543 );
mand \mul_6_19/U$157 ( \545 , \541 , \544 );
mor \mul_6_19/U$155 ( \546 , \540 , \545 );
mand \mul_6_19/U$152 ( \547 , \537 , \546 );
mor \mul_6_19/U$150 ( \548 , \536 , \547 );
mand \mul_6_19/U$147 ( \549 , \533 , \548 );
mor \mul_6_19/U$145 ( \550 , \532 , \549 );
mand \mul_6_19/U$142 ( \551 , \529 , \550 );
mor \mul_6_19/U$140 ( \552 , \528 , \551 );
mand \mul_6_19/U$137 ( \553 , \525 , \552 );
mor \mul_6_19/U$135 ( \554 , \524 , \553 );
mand \mul_6_19/U$132 ( \555 , \521 , \554 );
mor \mul_6_19/U$130 ( \556 , \520 , \555 );
mand \mul_6_19/U$127 ( \557 , \517 , \556 );
mor \mul_6_19/U$125 ( \558 , \516 , \557 );
mand \mul_6_19/U$122 ( \559 , \513 , \558 );
mor \mul_6_19/U$120 ( \560 , \512 , \559 );
mand \mul_6_19/U$117 ( \561 , \509 , \560 );
mor \mul_6_19/U$115 ( \562 , \508 , \561 );
mand \mul_6_19/U$105 ( \563 , \109_A[9] , \165_B[8] );
mand \mul_6_19/U$61 ( \564 , \562 , \563 );
mxor \mul_6_19/U$62 ( \565 , \562 , \563 );
mxor \mul_6_19/U$116 ( \566 , \509 , \560 );
mand \mul_6_19/U$106 ( \567 , \115_A[8] , \165_B[8] );
mand \mul_6_19/U$66 ( \568 , \566 , \567 );
mxor \mul_6_19/U$67 ( \569 , \566 , \567 );
mxor \mul_6_19/U$121 ( \570 , \513 , \558 );
mand \mul_6_19/U$107 ( \571 , \121_A[7] , \165_B[8] );
mand \mul_6_19/U$71 ( \572 , \570 , \571 );
mxor \mul_6_19/U$72 ( \573 , \570 , \571 );
mxor \mul_6_19/U$126 ( \574 , \517 , \556 );
mand \mul_6_19/U$108 ( \575 , \127_A[6] , \165_B[8] );
mand \mul_6_19/U$76 ( \576 , \574 , \575 );
mxor \mul_6_19/U$77 ( \577 , \574 , \575 );
mxor \mul_6_19/U$131 ( \578 , \521 , \554 );
mand \mul_6_19/U$109 ( \579 , \133_A[5] , \165_B[8] );
mand \mul_6_19/U$81 ( \580 , \578 , \579 );
mxor \mul_6_19/U$82 ( \581 , \578 , \579 );
mxor \mul_6_19/U$136 ( \582 , \525 , \552 );
mand \mul_6_19/U$110 ( \583 , \139_A[4] , \165_B[8] );
mand \mul_6_19/U$86 ( \584 , \582 , \583 );
mxor \mul_6_19/U$87 ( \585 , \582 , \583 );
mxor \mul_6_19/U$141 ( \586 , \529 , \550 );
mand \mul_6_19/U$111 ( \587 , \145_A[3] , \165_B[8] );
mand \mul_6_19/U$91 ( \588 , \586 , \587 );
mxor \mul_6_19/U$92 ( \589 , \586 , \587 );
mxor \mul_6_19/U$146 ( \590 , \533 , \548 );
mand \mul_6_19/U$112 ( \591 , \151_A[2] , \165_B[8] );
mand \mul_6_19/U$96 ( \592 , \590 , \591 );
mxor \mul_6_19/U$97 ( \593 , \590 , \591 );
mxor \mul_6_19/U$151 ( \594 , \537 , \546 );
mand \mul_6_19/U$113 ( \595 , \157_A[1] , \165_B[8] );
mand \mul_6_19/U$101 ( \596 , \594 , \595 );
mxor \mul_6_19/U$102 ( \597 , \594 , \595 );
mxor \mul_6_19/U$156 ( \598 , \541 , \544 );
mand \mul_6_19/U$114 ( \599 , \163_A[0] , \165_B[8] );
mand \mul_6_19/U$103 ( \600 , \598 , \599 );
mand \mul_6_19/U$100 ( \601 , \597 , \600 );
mor \mul_6_19/U$98 ( \602 , \596 , \601 );
mand \mul_6_19/U$95 ( \603 , \593 , \602 );
mor \mul_6_19/U$93 ( \604 , \592 , \603 );
mand \mul_6_19/U$90 ( \605 , \589 , \604 );
mor \mul_6_19/U$88 ( \606 , \588 , \605 );
mand \mul_6_19/U$85 ( \607 , \585 , \606 );
mor \mul_6_19/U$83 ( \608 , \584 , \607 );
mand \mul_6_19/U$80 ( \609 , \581 , \608 );
mor \mul_6_19/U$78 ( \610 , \580 , \609 );
mand \mul_6_19/U$75 ( \611 , \577 , \610 );
mor \mul_6_19/U$73 ( \612 , \576 , \611 );
mand \mul_6_19/U$70 ( \613 , \573 , \612 );
mor \mul_6_19/U$68 ( \614 , \572 , \613 );
mand \mul_6_19/U$65 ( \615 , \569 , \614 );
mor \mul_6_19/U$63 ( \616 , \568 , \615 );
mand \mul_6_19/U$60 ( \617 , \565 , \616 );
mor \mul_6_19/U$58 ( \618 , \564 , \617 );
mand \mul_6_19/U$48 ( \619 , \109_A[9] , \164_B[9] );
mand \mul_6_19/U$4 ( \620 , \618 , \619 );
mxor \mul_6_19/U$5 ( \621 , \618 , \619 );
mxor \mul_6_19/U$59 ( \622 , \565 , \616 );
mand \mul_6_19/U$49 ( \623 , \115_A[8] , \164_B[9] );
mand \mul_6_19/U$9 ( \624 , \622 , \623 );
mxor \mul_6_19/U$10 ( \625 , \622 , \623 );
mxor \mul_6_19/U$64 ( \626 , \569 , \614 );
mand \mul_6_19/U$50 ( \627 , \121_A[7] , \164_B[9] );
mand \mul_6_19/U$14 ( \628 , \626 , \627 );
mxor \mul_6_19/U$15 ( \629 , \626 , \627 );
mxor \mul_6_19/U$69 ( \630 , \573 , \612 );
mand \mul_6_19/U$51 ( \631 , \127_A[6] , \164_B[9] );
mand \mul_6_19/U$19 ( \632 , \630 , \631 );
mxor \mul_6_19/U$20 ( \633 , \630 , \631 );
mxor \mul_6_19/U$74 ( \634 , \577 , \610 );
mand \mul_6_19/U$52 ( \635 , \133_A[5] , \164_B[9] );
mand \mul_6_19/U$24 ( \636 , \634 , \635 );
mxor \mul_6_19/U$25 ( \637 , \634 , \635 );
mxor \mul_6_19/U$79 ( \638 , \581 , \608 );
mand \mul_6_19/U$53 ( \639 , \139_A[4] , \164_B[9] );
mand \mul_6_19/U$29 ( \640 , \638 , \639 );
mxor \mul_6_19/U$30 ( \641 , \638 , \639 );
mxor \mul_6_19/U$84 ( \642 , \585 , \606 );
mand \mul_6_19/U$54 ( \643 , \145_A[3] , \164_B[9] );
mand \mul_6_19/U$34 ( \644 , \642 , \643 );
mxor \mul_6_19/U$35 ( \645 , \642 , \643 );
mxor \mul_6_19/U$89 ( \646 , \589 , \604 );
mand \mul_6_19/U$55 ( \647 , \151_A[2] , \164_B[9] );
mand \mul_6_19/U$39 ( \648 , \646 , \647 );
mxor \mul_6_19/U$40 ( \649 , \646 , \647 );
mxor \mul_6_19/U$94 ( \650 , \593 , \602 );
mand \mul_6_19/U$56 ( \651 , \157_A[1] , \164_B[9] );
mand \mul_6_19/U$44 ( \652 , \650 , \651 );
mxor \mul_6_19/U$45 ( \653 , \650 , \651 );
mxor \mul_6_19/U$99 ( \654 , \597 , \600 );
mand \mul_6_19/U$57 ( \655 , \163_A[0] , \164_B[9] );
mand \mul_6_19/U$46 ( \656 , \654 , \655 );
mand \mul_6_19/U$43 ( \657 , \653 , \656 );
mor \mul_6_19/U$41 ( \658 , \652 , \657 );
mand \mul_6_19/U$38 ( \659 , \649 , \658 );
mor \mul_6_19/U$36 ( \660 , \648 , \659 );
mand \mul_6_19/U$33 ( \661 , \645 , \660 );
mor \mul_6_19/U$31 ( \662 , \644 , \661 );
mand \mul_6_19/U$28 ( \663 , \641 , \662 );
mor \mul_6_19/U$26 ( \664 , \640 , \663 );
mand \mul_6_19/U$23 ( \665 , \637 , \664 );
mor \mul_6_19/U$21 ( \666 , \636 , \665 );
mand \mul_6_19/U$18 ( \667 , \633 , \666 );
mor \mul_6_19/U$16 ( \668 , \632 , \667 );
mand \mul_6_19/U$13 ( \669 , \629 , \668 );
mor \mul_6_19/U$11 ( \670 , \628 , \669 );
mand \mul_6_19/U$8 ( \671 , \625 , \670 );
mor \mul_6_19/U$6 ( \672 , \624 , \671 );
mand \mul_6_19/U$3 ( \673 , \621 , \672 );
mor \mul_6_19/U$1 ( \674 , \620 , \673 );
mbuf \mul_6_19/Z[19] ( \675_Z[19] , \674 );
mxor \mul_6_19/U$2 ( \676 , \621 , \672 );
mbuf \mul_6_19/Z[18] ( \677_Z[18] , \676 );
mxor \mul_6_19/U$7 ( \678 , \625 , \670 );
mbuf \mul_6_19/Z[17] ( \679_Z[17] , \678 );
mxor \mul_6_19/U$12 ( \680 , \629 , \668 );
mbuf \mul_6_19/Z[16] ( \681_Z[16] , \680 );
mxor \mul_6_19/U$17 ( \682 , \633 , \666 );
mbuf \mul_6_19/Z[15] ( \683_Z[15] , \682 );
mxor \mul_6_19/U$22 ( \684 , \637 , \664 );
mbuf \mul_6_19/Z[14] ( \685_Z[14] , \684 );
mxor \mul_6_19/U$27 ( \686 , \641 , \662 );
mbuf \mul_6_19/Z[13] ( \687_Z[13] , \686 );
mxor \mul_6_19/U$32 ( \688 , \645 , \660 );
mbuf \mul_6_19/Z[12] ( \689_Z[12] , \688 );
mxor \mul_6_19/U$37 ( \690 , \649 , \658 );
mbuf \mul_6_19/Z[11] ( \691_Z[11] , \690 );
mxor \mul_6_19/U$42 ( \692 , \653 , \656 );
mbuf \mul_6_19/Z[10] ( \693_Z[10] , \692 );
mxor \mul_6_19/U$47 ( \694 , \654 , \655 );
mbuf \mul_6_19/Z[9] ( \695_Z[9] , \694 );
mxor \mul_6_19/U$104 ( \696 , \598 , \599 );
mbuf \mul_6_19/Z[8] ( \697_Z[8] , \696 );
mxor \mul_6_19/U$161 ( \698 , \542 , \543 );
mbuf \mul_6_19/Z[7] ( \699_Z[7] , \698 );
mxor \mul_6_19/U$218 ( \700 , \486 , \487 );
mbuf \mul_6_19/Z[6] ( \701_Z[6] , \700 );
mxor \mul_6_19/U$275 ( \702 , \430 , \431 );
mbuf \mul_6_19/Z[5] ( \703_Z[5] , \702 );
mxor \mul_6_19/U$332 ( \704 , \374 , \375 );
mbuf \mul_6_19/Z[4] ( \705_Z[4] , \704 );
mxor \mul_6_19/U$389 ( \706 , \318 , \319 );
mbuf \mul_6_19/Z[3] ( \707_Z[3] , \706 );
mxor \mul_6_19/U$446 ( \708 , \262 , \263 );
mbuf \mul_6_19/Z[2] ( \709_Z[2] , \708 );
mxor \mul_6_19/U$500 ( \710 , \207 , \208 );
mbuf \mul_6_19/Z[1] ( \711_Z[1] , \710 );
mand \mul_6_19/U$520 ( \712 , \163_A[0] , \173_B[0] );
mbuf \mul_6_19/Z[0] ( \713_Z[0] , \712 );
endmodule


//
// Conformal-LEC Version 19.20-d218 (25-Feb-2020)
//
module top( C, D, O);
input [1:0] C, D;
output [1:0] O;


m_DC \n6_5[1] ( O, C, D);

endmodule


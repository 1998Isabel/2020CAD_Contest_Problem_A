//
// Conformal-LEC Version 19.20-d218 (25-Feb-2020)
//
module top(\A[0][9] ,\A[0][8] ,\A[0][7] ,\A[0][6] ,\A[0][5] ,\A[0][4] ,\A[0][3] ,\A[0][2] ,\A[0][1] ,
        \A[0][0] ,\A[1][9] ,\A[1][8] ,\A[1][7] ,\A[1][6] ,\A[1][5] ,\A[1][4] ,\A[1][3] ,\A[1][2] ,\A[1][1] ,
        \A[1][0] ,\A[2][9] ,\A[2][8] ,\A[2][7] ,\A[2][6] ,\A[2][5] ,\A[2][4] ,\A[2][3] ,\A[2][2] ,\A[2][1] ,
        \A[2][0] ,\B[9] ,\B[8] ,\B[7] ,\B[6] ,\B[5] ,\B[4] ,\B[3] ,\B[2] ,\B[1] ,
        \B[0] ,\I[7] ,\I[6] ,\I[5] ,\I[4] ,\I[3] ,\I[2] ,\I[1] ,\I[0] ,\O[19] ,
        \O[18] ,\O[17] ,\O[16] ,\O[15] ,\O[14] ,\O[13] ,\O[12] ,\O[11] ,\O[10] ,\O[9] ,
        \O[8] ,\O[7] ,\O[6] ,\O[5] ,\O[4] ,\O[3] ,\O[2] ,\O[1] ,\O[0] );
input [1:0] \A[0][9] ,\A[0][8] ,\A[0][7] ,\A[0][6] ,\A[0][5] ,\A[0][4] ,\A[0][3] ,\A[0][2] ,\A[0][1] ,        \A[0][0] ,\A[1][9] ,\A[1][8] ,\A[1][7] ,\A[1][6] ,\A[1][5] ,\A[1][4] ,\A[1][3] ,\A[1][2] ,\A[1][1] ,        \A[1][0] ,\A[2][9] ,\A[2][8] ,\A[2][7] ,\A[2][6] ,\A[2][5] ,\A[2][4] ,\A[2][3] ,\A[2][2] ,\A[2][1] ,        \A[2][0] ,\B[9] ,\B[8] ,\B[7] ,\B[6] ,\B[5] ,\B[4] ,\B[3] ,\B[2] ,\B[1] ,        \B[0] ,\I[7] ,\I[6] ,\I[5] ,\I[4] ,\I[3] ,\I[2] ,\I[1] ,\I[0] ;
output [1:0] \O[19] ,\O[18] ,\O[17] ,\O[16] ,\O[15] ,\O[14] ,\O[13] ,\O[12] ,\O[11] ,        \O[10] ,\O[9] ,\O[8] ,\O[7] ,\O[6] ,\O[5] ,\O[4] ,\O[3] ,\O[2] ,\O[1] ,        \O[0] ;

wire [1:0] \69_ZERO , \70 , \71_ONE , \72 , \73 , \74 , \75 , \76 , \77 ,         \78 , \79 , \80 , \81 , \82 , \83 , \84 , \85 , \86 , \87 ,         \88 , \89 , \90 , \91 , \92 , \93 , \94 , \95 , \96 , \97 ,         \98 , \99 , \100 , \101 , \102 , \103 , \104 , \105 , \106 , \107 ,         \108 , \109 , \110 , \111 , \112 , \113 , \114 , \115 , \116 , \117 ,         \118 , \119 , \120 , \121 , \122 , \123 , \124 , \125 , \126 , \127 ,         \128 , \129 , \130 , \131 , \132 , \133 , \134 , \135 , \136 , \137 ,         \138 , \139 , \140 , \141 , \142 , \143 , \144 , \145 , \146 , \147 ,         \148 , \149 , \150 , \151 , \152 , \153 , \154 , \155 , \156 , \157 ,         \158 , \159 , \160 , \161 , \162 , \163 , \164 , \165 , \166 , \167 ,         \168 , \169 , \170 , \171 , \172 , \173 , \174 , \175 , \176 , \177 ,         \178 , \179 , \180 , \181 , \182 , \183 , \184 , \185 , \186 , \187 ,         \188 , \189 , \190 , \191 , \192 , \193 , \194 , \195 , \196 , \197 ,         \198 , \199 , \200 , \201 , \202 , \203 , \204 , \205 , \206 , \207 ,         \208 , \209 , \210 , \211 , \212 , \213 , \214 , \215 , \216 , \217 ,         \218 , \219 , \220 , \221 , \222 , \223 , \224 , \225 , \226 , \227 ,         \228 , \229 , \230 , \231 , \232 , \233 , \234 , \235 , \236 , \237 ,         \238 , \239 , \240 , \241 , \242 , \243 , \244 , \245 , \246 , \247 ,         \248 , \249 , \250 , \251 , \252 , \253 , \254 , \255 , \256 , \257 ,         \258 , \259 , \260 , \261 , \262 , \263 , \264 , \265 , \266 , \267 ,         \268 , \269 , \270 , \271 , \272 , \273 , \274 , \275 , \276 , \277 ,         \278 , \279 , \280 , \281 , \282 , \283 , \284 , \285 , \286 , \287 ,         \288 , \289 , \290 , \291 , \292 , \293 , \294 , \295 , \296 , \297 ,         \298 , \299 , \300 , \301 , \302 , \303 , \304 , \305 , \306 , \307 ,         \308 , \309 , \310 , \311 , \312 , \313 , \314 , \315 , \316 , \317 ,         \318 , \319 , \320 , \321 , \322 , \323 , \324 , \325 , \326 , \327 ,         \328 , \329 , \330 , \331 , \332 , \333 , \334 , \335 , \336 , \337 ,         \338 , \339 , \340 , \341 , \342 , \343 , \344 , \345 , \346 , \347 ,         \348 , \349 , \350 , \351 , \352 , \353 , \354 , \355 , \356 , \357 ,         \358 , \359 , \360 , \361 , \362 , \363 , \364 , \365 , \366 , \367 ,         \368 , \369 , \370 , \371 , \372 , \373 , \374 , \375 , \376 , \377 ,         \378 , \379 , \380 , \381 , \382 , \383 , \384 , \385 , \386 , \387 ,         \388 , \389 , \390 , \391 , \392 , \393 , \394 , \395 , \396 , \397 ,         \398 , \399 , \400 , \401 , \402 , \403 , \404 , \405 , \406 , \407 ,         \408 , \409 , \410 , \411 , \412 , \413 , \414 , \415 , \416 , \417 ,         \418 , \419 , \420 , \421 , \422 , \423 , \424 , \425 , \426 , \427 ,         \428 , \429 , \430 , \431 , \432 , \433 , \434 , \435 , \436 , \437 ,         \438 , \439 , \440 , \441 , \442 , \443 , \444 , \445 , \446 , \447 ,         \448 , \449 , \450 , \451 , \452 , \453 , \454 , \455 , \456 , \457 ,         \458 , \459 , \460 , \461 , \462 , \463 , \464 , \465 , \466 , \467 ,         \468 , \469 , \470 , \471 , \472 , \473 , \474 , \475 , \476 , \477 ,         \478 , \479 , \480 , \481 , \482 , \483 , \484 , \485 , \486 , \487 ,         \488 , \489 , \490 , \491 , \492 , \493 , \494 , \495 , \496 , \497 ,         \498 , \499 , \500 , \501 , \502 , \503 , \504 , \505 , \506 , \507 ,         \508 , \509 , \510 , \511 , \512 , \513 , \514 , \515 , \516 , \517 ,         \518 , \519 , \520 , \521 , \522 , \523 , \524 , \525 , \526 , \527 ,         \528 , \529 , \530 , \531 , \532 , \533 , \534 , \535 , \536 , \537 ,         \538 , \539 , \540 , \541 , \542 , \543 , \544 , \545 , \546 , \547 ,         \548 , \549 , \550 , \551 , \552 , \553 , \554 , \555 , \556 , \557 ,         \558 , \559 , \560 , \561 , \562 , \563 , \564 , \565 , \566 , \567 ,         \568 , \569 , \570 , \571 , \572 , \573 , \574 , \575 , \576 , \577 ,         \578 , \579 , \580 , \581 , \582 , \583 , \584 , \585 , \586 , \587 ,         \588 , \589 , \590 , \591 , \592 , \593 , \594 , \595 , \596 , \597 ,         \598 , \599 , \600 , \601 , \602 , \603 , \604 , \605 , \606 , \607 ,         \608 , \609 , \610 , \611 , \612 , \613 , \614 , \615 , \616 , \617 ,         \618 , \619 , \620 , \621 , \622 , \623 , \624 , \625 , \626 , \627 ,         \628 , \629 , \630 , \631 , \632 , \633 , \634 , \635 , \636 , \637 ,         \638 , \639 , \640 , \641 , \642 , \643 , \644 , \645 , \646 , \647 ,         \648 , \649 , \650 , \651 , \652 , \653 , \654 , \655 , \656 , \657 ,         \658 , \659 , \660 , \661 , \662 , \663 , \664 , \665 , \666 , \667 ,         \668 , \669 , \670 , \671 , \672 , \673 , \674 , \675 , \676 , \677 ,         \678 , \679 , \680 , \681 , \682 , \683 , \684 , \685 , \686 , \687 ,         \688 , \689 , \690 , \691 , \692 , \693 , \694 , \695 , \696 , \697 ,         \698 , \699 , \700 , \701 , \702 , \703 , \704 , \705 , \706 , \707 ,         \708 , \709 , \710 , \711 , \712 , \713 , \714 , \715 , \716 , \717 ,         \718 , \719 , \720 , \721 , \722 , \723 , \724 , \725 , \726 , \727 ,         \728 , \729 , \730 , \731 , \732 , \733 , \734 , \735 , \736 , \737 ,         \738 , \739 , \740 , \741 , \742 , \743 , \744 , \745 , \746 , \747 ,         \748 , \749 , \750 , \751 , \752 , \753 , \754 , \755 , \756 , \757 ,         \758 , \759 , \760 , \761 , \762 , \763 , \764 , \765 , \766 , \767 ,         \768 , \769 , \770 , \771 , \772 , \773 , \774 , \775 , \776 , \777 ,         \778 , \779 , \780 , \781 , \782 , \783 , \784 , \785 , \786 , \787 ,         \788 , \789 , \790 , \791 , \792 , \793 , \794 , \795 , \796 , \797 ,         \798 , \799 , \800 , \801 , \802 , \803 , \804 , \805 , \806 , \807 ,         \808 , \809 , \810 , \811 , \812 , \813 , \814 , \815 , \816 , \817 ,         \818 , \819 , \820 , \821 , \822 , \823 , \824 , \825 , \826 , \827 ,         \828 , \829 , \830 , \831 , \832 , \833 , \834 , \835 , \836 , \837 ,         \838 , \839 , \840 , \841 , \842 , \843 , \844 , \845 , \846 , \847 ,         \848 , \849 , \850 , \851 , \852 , \853 , \854 , \855 , \856 , \857 ,         \858 , \859 , \860 , \861 , \862 , \863 , \864 , \865 , \866 , \867 ,         \868 , \869 , \870 , \871 , \872 , \873 , \874 , \875 , \876 , \877 ,         \878 , \879 , \880 , \881 , \882 , \883 , \884 , \885 , \886 , \887 ,         \888 , \889 , \890 , \891 , \892 , \893 , \894 , \895 , \896 , \897 ,         \898 , \899 , \900 , \901 , \902 , \903 , \904 , \905 , \906 , \907 ,         \908 , \909 , \910 , \911 , \912 , \913 , \914 , \915 , \916 , \917 ,         \918 , \919 , \920 , \921 , \922 , \923 , \924 , \925 , \926 , \927 ,         \928 , \929 , \930 , \931 , \932 , \933 , \934 , \935 , \936 , \937 ,         \938 , \939 , \940 , \941 , \942 , \943 , \944 , \945 , \946 , \947 ,         \948 , \949 , \950 , \951 , \952 , \953 , \954 , \955 , \956 , \957 ,         \958 , \959 , \960 , \961 , \962 , \963 , \964 , \965 , \966 , \967 ,         \968 , \969 , \970 , \971 , \972 , \973 , \974 , \975 , \976 , \977 ,         \978 , \979 , \980 , \981 , \982 , \983 , \984 , \985 , \986 , \987 ,         \988 , \989 , \990 , \991 , \992 , \993 , \994 , \995 , \996 , \997 ,         \998 , \999 , \1000 , \1001 , \1002 , \1003 , \1004 , \1005 , \1006 , \1007 ,         \1008 , \1009 , \1010 , \1011 , \1012 , \1013 , \1014 , \1015 , \1016 , \1017 ,         \1018 , \1019 , \1020 , \1021 , \1022 , \1023 , \1024 , \1025 , \1026 , \1027 ,         \1028 , \1029 , \1030 , \1031 , \1032 , \1033 , \1034 , \1035 , \1036 , \1037 ,         \1038 , \1039 , \1040 , \1041 , \1042 , \1043 , \1044 , \1045 , \1046 , \1047 ,         \1048 , \1049 , \1050 , \1051 , \1052 , \1053 , \1054 , \1055 , \1056 , \1057 ,         \1058 , \1059 , \1060 , \1061 , \1062 , \1063 , \1064 , \1065 , \1066 , \1067 ,         \1068 , \1069 , \1070 , \1071 , \1072 , \1073 , \1074 , \1075 ;
mbuf \U$labaj121 ( \O[19] , \943 );
mbuf \U$labaj122 ( \O[18] , \949 );
mbuf \U$labaj123 ( \O[17] , \969 );
mbuf \U$labaj124 ( \O[16] , \1073 );
mbuf \U$labaj125 ( \O[15] , \985 );
mbuf \U$labaj126 ( \O[14] , \1074 );
mbuf \U$labaj127 ( \O[13] , \997 );
mbuf \U$labaj128 ( \O[12] , \1075 );
mbuf \U$labaj129 ( \O[11] , \1010 );
mbuf \U$labaj130 ( \O[10] , \1017 );
mbuf \U$labaj131 ( \O[9] , \1024 );
mbuf \U$labaj132 ( \O[8] , \1030 );
mbuf \U$labaj133 ( \O[7] , \1039 );
mbuf \U$labaj134 ( \O[6] , \1047 );
mbuf \U$labaj135 ( \O[5] , \1053 );
mbuf \U$labaj136 ( \O[4] , \1059 );
mbuf \U$labaj137 ( \O[3] , \1065 );
mbuf \U$labaj138 ( \O[2] , \1067 );
mbuf \U$labaj139 ( \O[1] , \1071 );
mbuf \U$labaj140 ( \O[0] , \1072 );
mnot \g11877/U$3 ( \72 , \A[0][5] );
mnor \g3/U$1 ( \73 , \I[1] , \I[0] );
mnot \g11877/U$4 ( \74 , \73 );
mor \g11877/U$2 ( \75 , \72 , \74 );
mand \g707/U$2 ( \76 , \A[1][5] , \I[0] );
mand \g707/U$3 ( \77 , \A[2][5] , \I[1] );
mnor \g707/U$1 ( \78 , \76 , \77 );
mnand \g11877/U$1 ( \79 , \75 , \78 );
mbuf \g678/U$1 ( \80 , \79 );
mnand \mul_6_19_g11737/U$1 ( \81 , \80 , \B[9] );
mnot \g11989/U$2 ( \82 , \A[0][7] );
mnor \g11989/U$1 ( \83 , \82 , \I[0] , \I[1] );
mnand \g723/U$1 ( \84 , \A[2][7] , \I[1] );
mnand \g724/U$1 ( \85 , \A[1][7] , \I[0] );
mnand \g709/U$1 ( \86 , \84 , \85 );
mnor \g677/U$1 ( \87 , \83 , \86 );
mnot \g676/U$1 ( \88 , \87 );
mnand \mul_6_19_g11747/U$1 ( \89 , \88 , \B[7] );
mxor \mul_6_19_g11474/U$4 ( \90 , \81 , \89 );
mnand \mul_6_19_g11709/U$1 ( \91 , \80 , \B[8] );
mnor \g11968/U$1 ( \92 , \I[1] , \I[0] );
mnot \g12005/U$3 ( \93 , \92 );
mnot \g12005/U$4 ( \94 , \A[0][4] );
mor \g12005/U$2 ( \95 , \93 , \94 );
mand \g711/U$2 ( \96 , \A[1][4] , \I[0] );
mand \g711/U$3 ( \97 , \A[2][4] , \I[1] );
mnor \g711/U$1 ( \98 , \96 , \97 );
mnand \g12005/U$1 ( \99 , \95 , \98 );
mbuf \g687/U$1 ( \100 , \99 );
mnand \mul_6_19_g11868/U$1 ( \101 , \100 , \B[9] );
mxor \mul_6_19_g11512/U$4 ( \102 , \91 , \101 );
mnand \mul_6_19_g11742/U$1 ( \103 , \88 , \B[6] );
mand \mul_6_19_g11512/U$3 ( \104 , \102 , \103 );
mand \mul_6_19_g11512/U$5 ( \105 , \91 , \101 );
mor \mul_6_19_g11512/U$2 ( \106 , \104 , \105 );
mand \mul_6_19_g11474/U$3 ( \107 , \90 , \106 );
mand \mul_6_19_g11474/U$5 ( \108 , \81 , \89 );
mor \mul_6_19_g11474/U$2 ( \109 , \107 , \108 );
mnand \mul_6_19_g11633/U$1 ( \110 , \88 , \B[8] );
mnor \g11970/U$1 ( \111 , \I[1] , \I[0] );
mnot \g12006/U$3 ( \112 , \111 );
mnot \g12006/U$4 ( \113 , \A[0][6] );
mor \g12006/U$2 ( \114 , \112 , \113 );
mand \g703/U$2 ( \115 , \A[1][6] , \I[0] );
mand \g703/U$3 ( \116 , \A[2][6] , \I[1] );
mnor \g703/U$1 ( \117 , \115 , \116 );
mnand \g12006/U$1 ( \118 , \114 , \117 );
mbuf \g689/U$1 ( \119 , \118 );
mnand \mul_6_19_g11672/U$1 ( \120 , \119 , \B[8] );
mnor \g11962/U$1 ( \121 , \I[1] , \I[0] );
mnot \g12001/U$3 ( \122 , \121 );
mnot \g12001/U$4 ( \123 , \A[0][9] );
mor \g12001/U$2 ( \124 , \122 , \123 );
mand \g710/U$2 ( \125 , \A[1][9] , \I[0] );
mand \g710/U$3 ( \126 , \A[2][9] , \I[1] );
mnor \g710/U$1 ( \127 , \125 , \126 );
mnand \g12001/U$1 ( \128 , \124 , \127 );
mbuf \g674/U$1 ( \129 , \128 );
mnand \mul_6_19_g11636/U$1 ( \130 , \129 , \B[5] );
mxor \mul_6_19_g11513/U$4 ( \131 , \120 , \130 );
mnor \g11966/U$1 ( \132 , \I[1] , \I[0] );
mnot \g12004/U$3 ( \133 , \132 );
mnot \g12004/U$4 ( \134 , \A[0][8] );
mor \g12004/U$2 ( \135 , \133 , \134 );
mand \g705/U$2 ( \136 , \A[1][8] , \I[0] );
mand \g705/U$3 ( \137 , \A[2][8] , \I[1] );
mnor \g705/U$1 ( \138 , \136 , \137 );
mnand \g12004/U$1 ( \139 , \135 , \138 );
mbuf \mul_6_19_g11756/U$1 ( \140 , \139 );
mnand \mul_6_19_g11685/U$1 ( \141 , \140 , \B[6] );
mand \mul_6_19_g11513/U$3 ( \142 , \131 , \141 );
mand \mul_6_19_g11513/U$5 ( \143 , \120 , \130 );
mor \mul_6_19_g11513/U$2 ( \144 , \142 , \143 );
mxor \mul_6_19_g11440/U$1 ( \145 , \110 , \144 );
mnand \mul_6_19_g11749/U$1 ( \146 , \140 , \B[7] );
mnand \mul_6_19_g11637/U$1 ( \147 , \129 , \B[6] );
mxor \mul_6_19_g11530/U$1 ( \148 , \146 , \147 );
mnand \mul_6_19_g11719/U$1 ( \149 , \119 , \B[9] );
mxor \mul_6_19_g11530/U$1_r1 ( \150 , \148 , \149 );
mxor \mul_6_19_g11440/U$1_r1 ( \151 , \145 , \150 );
mxor \mul_6_19_g11371/U$1 ( \152 , \109 , \151 );
mxor \mul_6_19_g11474/U$1 ( \153 , \81 , \89 );
mxor \mul_6_19_g11474/U$1_r1 ( \154 , \153 , \106 );
mxor \mul_6_19_g11513/U$1 ( \155 , \120 , \130 );
mxor \mul_6_19_g11513/U$1_r1 ( \156 , \155 , \141 );
mnand \mul_6_19_g11450/U$1 ( \157 , \154 , \156 );
mnand \mul_6_19_g11720/U$1 ( \158 , \140 , \B[5] );
mnand \mul_6_19_g11686/U$1 ( \159 , \129 , \B[4] );
mxor \mul_6_19_g11516/U$4 ( \160 , \158 , \159 );
mnand \mul_6_19_g11625/U$1 ( \161 , \119 , \B[7] );
mand \mul_6_19_g11516/U$3 ( \162 , \160 , \161 );
mand \mul_6_19_g11516/U$5 ( \163 , \158 , \159 );
mor \mul_6_19_g11516/U$2 ( \164 , \162 , \163 );
mnot \mul_6_19_g11515/U$1 ( \165 , \164 );
mand \mul_6_19_g11425/U$2 ( \166 , \157 , \165 );
mnor \mul_6_19_g11455/U$1 ( \167 , \154 , \156 );
mnor \mul_6_19_g11425/U$1 ( \168 , \166 , \167 );
mxor \mul_6_19_g11371/U$1_r1 ( \169 , \152 , \168 );
mnot \mul_6_19_g11768/U$2 ( \170 , \169 );
mxor \mul_6_19_g11516/U$1 ( \171 , \158 , \159 );
mxor \mul_6_19_g11516/U$1_r1 ( \172 , \171 , \161 );
mnand \mul_6_19_g11715/U$1 ( \173 , \139 , \B[4] );
mnot \mul_6_19_g11561/U$3 ( \174 , \173 );
mnand \mul_6_19_g11985/U$1 ( \175 , \129 , \B[3] );
mnot \mul_6_19_g11561/U$4 ( \176 , \175 );
mor \mul_6_19_g11561/U$2 ( \177 , \174 , \176 );
mand \mul_6_19_g11689/U$1 ( \178 , \119 , \B[6] );
mnand \mul_6_19_g11561/U$1 ( \179 , \177 , \178 );
mnot \mul_6_19_g11602/U$2 ( \180 , \175 );
mnot \mul_6_19_g11714/U$1 ( \181 , \173 );
mnand \mul_6_19_g11602/U$1 ( \182 , \180 , \181 );
mnand \mul_6_19_g11533/U$1 ( \183 , \179 , \182 );
mnot \mul_6_19_g11528/U$1 ( \184 , \183 );
mnand \mul_6_19_g11497/U$1 ( \185 , \172 , \184 );
mnot \mul_6_19_g2/U$3 ( \186 , \185 );
mnand \mul_6_19_g11660/U$1 ( \187 , \80 , \B[7] );
mnand \mul_6_19_g11630/U$1 ( \188 , \88 , \B[5] );
mand \g11982/U$1 ( \189 , \187 , \188 );
mnand \mul_6_19_g11676/U$1 ( \190 , \100 , \B[8] );
mor \g11981/U$2 ( \191 , \189 , \190 );
mor \mul_6_19_g11784/U$1 ( \192 , \188 , \187 );
mnand \g11981/U$1 ( \193 , \191 , \192 );
mnot \mul_6_19_g2/U$4 ( \194 , \193 );
mor \mul_6_19_g2/U$2 ( \195 , \186 , \194 );
mor \mul_6_19_g2/U$5 ( \196 , \172 , \184 );
mnand \mul_6_19_g2/U$1 ( \197 , \195 , \196 );
mand \mul_6_19_g11493/U$2 ( \198 , \156 , \164 );
mnot \mul_6_19_g11493/U$4 ( \199 , \156 );
mand \mul_6_19_g11493/U$3 ( \200 , \199 , \165 );
mnor \mul_6_19_g11493/U$1 ( \201 , \198 , \200 );
mand \mul_6_19_g11449/U$2 ( \202 , \201 , \154 );
mnot \mul_6_19_g11449/U$4 ( \203 , \201 );
mnot \fopt11848/U$1 ( \204 , \154 );
mand \mul_6_19_g11449/U$3 ( \205 , \203 , \204 );
mor \mul_6_19_g11449/U$1 ( \206 , \202 , \205 );
mxor \mul_6_19_g11355/U$4 ( \207 , \197 , \206 );
mxor \mul_6_19_g11512/U$1 ( \208 , \91 , \101 );
mxor \mul_6_19_g11512/U$1_r1 ( \209 , \208 , \103 );
mnot \mul_6_19_g11415/U$3 ( \210 , \209 );
mnot \mul_6_19_g11526/U$1 ( \211 , \183 );
mnot \mul_6_19_g11492/U$3 ( \212 , \211 );
mnot \mul_6_19_g11492/U$4 ( \213 , \193 );
mand \mul_6_19_g11492/U$2 ( \214 , \212 , \213 );
mand \mul_6_19_g11492/U$5 ( \215 , \193 , \184 );
mnor \mul_6_19_g11492/U$1 ( \216 , \214 , \215 );
mnot \mul_6_19_g11467/U$3 ( \217 , \216 );
mnot \mul_6_19_g11514/U$1 ( \218 , \172 );
mnot \mul_6_19_g11467/U$4 ( \219 , \218 );
mor \mul_6_19_g11467/U$2 ( \220 , \217 , \219 );
mnot \mul_6_19_g11775/U$2 ( \221 , \216 );
mnand \mul_6_19_g11775/U$1 ( \222 , \221 , \172 );
mnand \mul_6_19_g11467/U$1 ( \223 , \220 , \222 );
mnot \mul_6_19_g11442/U$1 ( \224 , \223 );
mnot \mul_6_19_g11415/U$4 ( \225 , \224 );
mor \mul_6_19_g11415/U$2 ( \226 , \210 , \225 );
mnot \g735/U$1 ( \227 , \A[0][3] );
mnor \g701/U$1 ( \228 , \227 , \I[0] , \I[1] );
mnand \g715/U$1 ( \229 , \A[2][3] , \I[1] );
mnand \g714/U$1 ( \230 , \A[1][3] , \I[0] );
mnand \g712/U$1 ( \231 , \229 , \230 );
mnor \g692/U$1 ( \232 , \228 , \231 );
mnot \g691/U$1 ( \233 , \232 );
mbuf \mul_6_19_g11754/U$1 ( \234 , \233 );
mnand \mul_6_19_g11727/U$1 ( \235 , \234 , \B[9] );
mnand \mul_6_19_g11674/U$1 ( \236 , \139 , \B[3] );
mnand \mul_6_19_g11935/U$1 ( \237 , \119 , \B[5] );
mxor \mul_6_19_g11510/U$4 ( \238 , \236 , \237 );
mnand \mul_6_19_g11701/U$1 ( \239 , \129 , \B[2] );
mand \mul_6_19_g11510/U$3 ( \240 , \238 , \239 );
mand \mul_6_19_g11510/U$5 ( \241 , \236 , \237 );
mor \mul_6_19_g11510/U$2 ( \242 , \240 , \241 );
mxor \mul_6_19_g11439/U$4 ( \243 , \235 , \242 );
mnand \mul_6_19_g11635/U$1 ( \244 , \80 , \B[6] );
mnor \g11960/U$1 ( \245 , \I[1] , \I[0] );
mnot \g12002/U$3 ( \246 , \245 );
mnot \g12002/U$4 ( \247 , \A[0][2] );
mor \g12002/U$2 ( \248 , \246 , \247 );
mand \g704/U$2 ( \249 , \A[1][2] , \I[0] );
mand \g704/U$3 ( \250 , \A[2][2] , \I[1] );
mnor \g704/U$1 ( \251 , \249 , \250 );
mnand \g12002/U$1 ( \252 , \248 , \251 );
mbuf \g680/U$1 ( \253 , \252 );
mnand \mul_6_19_g11744/U$1 ( \254 , \253 , \B[9] );
mxor \mul_6_19_g11532/U$4 ( \255 , \244 , \254 );
mnand \mul_6_19_g11751/U$1 ( \256 , \88 , \B[4] );
mand \mul_6_19_g11532/U$3 ( \257 , \255 , \256 );
mand \mul_6_19_g11532/U$5 ( \258 , \244 , \254 );
mor \mul_6_19_g11532/U$2 ( \259 , \257 , \258 );
mand \mul_6_19_g11439/U$3 ( \260 , \243 , \259 );
mand \mul_6_19_g11439/U$5 ( \261 , \235 , \242 );
mor \mul_6_19_g11439/U$2 ( \262 , \260 , \261 );
mnot \mul_6_19_g11438/U$1 ( \263 , \262 );
mnand \mul_6_19_g11415/U$1 ( \264 , \226 , \263 );
mnot \mul_6_19_g11420/U$2 ( \265 , \209 );
mnand \mul_6_19_g11420/U$1 ( \266 , \265 , \223 );
mnand \mul_6_19_g11404/U$1 ( \267 , \264 , \266 );
mand \mul_6_19_g11355/U$3 ( \268 , \207 , \267 );
mand \mul_6_19_g11355/U$5 ( \269 , \197 , \206 );
mor \mul_6_19_g11355/U$2 ( \270 , \268 , \269 );
mnor \mul_6_19_g11768/U$1 ( \271 , \170 , \270 );
mnot \fopt11898/U$1 ( \272 , \271 );
mnot \g11950/U$2 ( \273 , \272 );
mnot \mul_6_19_g11766/U$2 ( \274 , \270 );
mnor \mul_6_19_g11766/U$1 ( \275 , \274 , \169 );
mnor \g11950/U$1 ( \276 , \273 , \275 );
mnot \mul_6_19_g11329/U$1 ( \277 , \276 );
mor \U$5 ( \278 , \I[7] , \I[6] , \I[5] , \I[4] , \I[3] , \I[2] , \I[1] , \I[0] );
mand \U$4 ( \279 , \B[9] , \B[8] , \B[7] , \B[6] , \B[5] , \B[4] , \B[3] , \B[2] , \B[1] , \B[0] );
mnot \U$3 ( \280 , \279 );
mor \U$2 ( \281 , \278 , \280 );
m_HMUX \U$1 ( \282 , 1'b1 , \277 , \281 );
mnot \g11939/U$2 ( \283 , \A[0][1] );
mnor \g11939/U$1 ( \284 , \283 , \I[0] , \I[1] );
mnand \g718/U$1 ( \285 , \A[2][1] , \I[1] );
mnand \g720/U$1 ( \286 , \A[1][1] , \I[0] );
mnand \g706/U$1 ( \287 , \285 , \286 );
mnor \g683/U$1 ( \288 , \284 , \287 );
mnot \g682/U$1 ( \289 , \288 );
mnor \g11964/U$1 ( \290 , \I[1] , \I[0] );
mnand \g11963/U$1 ( \291 , \290 , \A[0][0] );
mand \g708/U$2 ( \292 , \A[1][0] , \I[0] );
mand \g708/U$3 ( \293 , \A[2][0] , \I[1] );
mnor \g708/U$1 ( \294 , \292 , \293 );
mnand \g685/U$1 ( \295 , \291 , \294 );
mbuf \g684/U$1 ( \296 , \295 );
mnand \mul_6_19_g11706/U$1 ( \297 , \129 , \B[8] );
mnand \mul_6_19_g11621/U$1 ( \298 , \140 , \B[9] );
mxor \mul_6_19_g11476/U$4 ( \299 , \297 , \298 );
mnand \mul_6_19_g11687/U$1 ( \300 , \129 , \B[7] );
mnand \mul_6_19_g11634/U$1 ( \301 , \88 , \B[9] );
mxor \mul_6_19_g11520/U$4 ( \302 , \300 , \301 );
mnand \mul_6_19_g11667/U$1 ( \303 , \140 , \B[8] );
mand \mul_6_19_g11520/U$3 ( \304 , \302 , \303 );
mand \mul_6_19_g11520/U$5 ( \305 , \300 , \301 );
mor \mul_6_19_g11520/U$2 ( \306 , \304 , \305 );
mand \mul_6_19_g11476/U$3 ( \307 , \299 , \306 );
mand \mul_6_19_g11476/U$5 ( \308 , \297 , \298 );
mor \mul_6_19_g11476/U$2 ( \309 , \307 , \308 );
mnand \mul_6_19_g11753/U$1 ( \310 , \129 , \B[9] );
mnand \mul_6_19_g11454/U$1 ( \311 , \309 , \310 );
mnot \mul_6_19_g11245/U$3 ( \312 , \311 );
mxor \mul_6_19_g11986/U$1 ( \313 , \187 , \190 );
mxor \mul_6_19_g11986/U$1_r1 ( \314 , \313 , \188 );
mxor \g11956/U$1 ( \315 , \175 , \173 );
mxnor \g11956/U$1_r1 ( \316 , \315 , \178 );
mand \mul_6_19_g11456/U$2 ( \317 , \314 , \316 );
mnand \mul_6_19_g11662/U$1 ( \318 , \233 , \B[8] );
mnand \mul_6_19_g11869/U$1 ( \319 , \100 , \B[7] );
mxor \mul_6_19_g11519/U$4 ( \320 , \318 , \319 );
mand \mul_6_19_g11703/U$1 ( \321 , \129 , \B[1] );
mand \mul_6_19_g11718/U$1 ( \322 , \139 , \B[2] );
mnand \mul_6_19_g11610/U$1 ( \323 , \321 , \322 );
mand \mul_6_19_g11519/U$3 ( \324 , \320 , \323 );
mand \mul_6_19_g11519/U$5 ( \325 , \318 , \319 );
mor \mul_6_19_g11519/U$2 ( \326 , \324 , \325 );
mnor \mul_6_19_g11456/U$1 ( \327 , \317 , \326 );
mnot \fopt11893/U$1 ( \328 , \316 );
mnot \mul_6_19_g11529/U$1 ( \329 , \314 );
mand \mul_6_19_g11475/U$2 ( \330 , \328 , \329 );
mnor \mul_6_19_g11433/U$1 ( \331 , \327 , \330 );
mnot \mul_6_19_g11340/U$3 ( \332 , \331 );
mxor \mul_6_19_g11402/U$1 ( \333 , \209 , \262 );
mxnor \mul_6_19_g11402/U$1_r1 ( \334 , \333 , \223 );
mnot \mul_6_19_g11340/U$4 ( \335 , \334 );
mor \mul_6_19_g11340/U$2 ( \336 , \332 , \335 );
mxor \mul_6_19_g11439/U$1 ( \337 , \235 , \242 );
mxor \mul_6_19_g11439/U$1_r1 ( \338 , \337 , \259 );
mxor \mul_6_19_g11510/U$1 ( \339 , \236 , \237 );
mxor \mul_6_19_g11510/U$1_r1 ( \340 , \339 , \239 );
mnot \g11949/U$2 ( \341 , \340 );
mnand \mul_6_19_g11717/U$1 ( \342 , \119 , \B[4] );
mnot \mul_6_19_g11560/U$3 ( \343 , \342 );
mnand \mul_6_19_g11934/U$1 ( \344 , \253 , \B[8] );
mnot \mul_6_19_g11560/U$4 ( \345 , \344 );
mor \mul_6_19_g11560/U$2 ( \346 , \343 , \345 );
mand \mul_6_19_g11693/U$1 ( \347 , \289 , \B[9] );
mnand \mul_6_19_g11560/U$1 ( \348 , \346 , \347 );
mnot \mul_6_19_g11788/U$2 ( \349 , \342 );
mnot \mul_6_19_g11734/U$1 ( \350 , \344 );
mnand \mul_6_19_g11788/U$1 ( \351 , \349 , \350 );
mnand \mul_6_19_g11534/U$1 ( \352 , \348 , \351 );
mnand \g11949/U$1 ( \353 , \341 , \352 );
mnot \mul_6_19_g11517/U$1 ( \354 , \352 );
mnot \mul_6_19_g11482/U$3 ( \355 , \354 );
mnot \mul_6_19_g11482/U$4 ( \356 , \340 );
mor \mul_6_19_g11482/U$2 ( \357 , \355 , \356 );
mnand \mul_6_19_g11650/U$1 ( \358 , \80 , \B[5] );
mnot \mul_6_19_g11562/U$3 ( \359 , \358 );
mnand \mul_6_19_g11632/U$1 ( \360 , \88 , \B[3] );
mnot \mul_6_19_g11562/U$4 ( \361 , \360 );
mor \mul_6_19_g11562/U$2 ( \362 , \359 , \361 );
mnand \mul_6_19_g11867/U$1 ( \363 , \100 , \B[6] );
mnot \mul_6_19_g11640/U$1 ( \364 , \363 );
mnand \mul_6_19_g11562/U$1 ( \365 , \362 , \364 );
mor \mul_6_19_g11781/U$1 ( \366 , \360 , \358 );
mnand \mul_6_19_g11535/U$1 ( \367 , \365 , \366 );
mnand \mul_6_19_g11482/U$1 ( \368 , \357 , \367 );
mand \g11936/U$1 ( \369 , \353 , \368 );
mxor \mul_6_19_g11394/U$4 ( \370 , \338 , \369 );
mxor \mul_6_19_g11532/U$1 ( \371 , \244 , \254 );
mxor \mul_6_19_g11532/U$1_r1 ( \372 , \371 , \256 );
mxor \mul_6_19_g11519/U$1 ( \373 , \318 , \319 );
mxor \mul_6_19_g11519/U$1_r1 ( \374 , \373 , \323 );
mxor \mul_6_19_g11430/U$4 ( \375 , \372 , \374 );
mnand \mul_6_19_g11694/U$1 ( \376 , \234 , \B[7] );
mnand \mul_6_19_g11721/U$1 ( \377 , \129 , \B[0] );
mnot \mul_6_19_g11606/U$2 ( \378 , \377 );
mand \mul_6_19_g11695/U$1 ( \379 , \139 , \B[1] );
mnand \mul_6_19_g11606/U$1 ( \380 , \378 , \379 );
mxor \mul_6_19_g11487/U$4 ( \381 , \376 , \380 );
mxnor \g11818/U$1 ( \382 , \322 , \321 );
mand \mul_6_19_g11487/U$3 ( \383 , \381 , \382 );
mand \mul_6_19_g11487/U$5 ( \384 , \376 , \380 );
mor \mul_6_19_g11487/U$2 ( \385 , \383 , \384 );
mand \mul_6_19_g11430/U$3 ( \386 , \375 , \385 );
mand \mul_6_19_g11430/U$5 ( \387 , \372 , \374 );
mor \mul_6_19_g11430/U$2 ( \388 , \386 , \387 );
mand \mul_6_19_g11394/U$3 ( \389 , \370 , \388 );
mand \mul_6_19_g11394/U$5 ( \390 , \338 , \369 );
mor \mul_6_19_g11394/U$2 ( \391 , \389 , \390 );
mnot \mul_6_19_g11393/U$1 ( \392 , \391 );
mnand \mul_6_19_g11340/U$1 ( \393 , \336 , \392 );
mor \g11944/U$1 ( \394 , \334 , \331 );
mnand \mul_6_19_g11332/U$1 ( \395 , \393 , \394 );
mxor \mul_6_19_g11355/U$1 ( \396 , \197 , \206 );
mxor \mul_6_19_g11355/U$1_r1 ( \397 , \396 , \267 );
mor \mul_6_19_g11764/U$1 ( \398 , \395 , \397 );
mnand \mul_6_19_g11858/U$1 ( \399 , \398 , \272 );
mxor \mul_6_19_g11530/U$4 ( \400 , \146 , \147 );
mand \mul_6_19_g11530/U$3 ( \401 , \400 , \149 );
mand \mul_6_19_g11530/U$5 ( \402 , \146 , \147 );
mor \mul_6_19_g11530/U$2 ( \403 , \401 , \402 );
mxor \mul_6_19_g11520/U$1 ( \404 , \300 , \301 );
mxor \mul_6_19_g11520/U$1_r1 ( \405 , \404 , \303 );
mxor \mul_6_19_g11407/U$4 ( \406 , \403 , \405 );
mxor \mul_6_19_g11440/U$4 ( \407 , \110 , \144 );
mand \mul_6_19_g11440/U$3 ( \408 , \407 , \150 );
mand \mul_6_19_g11440/U$5 ( \409 , \110 , \144 );
mor \mul_6_19_g11440/U$2 ( \410 , \408 , \409 );
mand \mul_6_19_g11407/U$3 ( \411 , \406 , \410 );
mand \mul_6_19_g11407/U$5 ( \412 , \403 , \405 );
mor \mul_6_19_g11407/U$2 ( \413 , \411 , \412 );
mxor \mul_6_19_g11476/U$1 ( \414 , \297 , \298 );
mxor \mul_6_19_g11476/U$1_r1 ( \415 , \414 , \306 );
mnand \mul_6_19_g11395/U$1 ( \416 , \413 , \415 );
mxor \mul_6_19_g11371/U$4 ( \417 , \109 , \151 );
mand \mul_6_19_g11371/U$3 ( \418 , \417 , \168 );
mand \mul_6_19_g11371/U$5 ( \419 , \109 , \151 );
mor \mul_6_19_g11371/U$2 ( \420 , \418 , \419 );
mxor \mul_6_19_g11407/U$1 ( \421 , \403 , \405 );
mxor \mul_6_19_g11407/U$1_r1 ( \422 , \421 , \410 );
mnand \mul_6_19_g11357/U$1 ( \423 , \420 , \422 );
mnand \mul_6_19_g11344/U$1 ( \424 , \416 , \423 );
mnor \mul_6_19_g11277/U$1 ( \425 , \399 , \424 );
mnot \mul_6_19_g11762/U$2 ( \426 , \425 );
mxor \mul_6_19_g11394/U$1 ( \427 , \338 , \369 );
mxor \mul_6_19_g11394/U$1_r1 ( \428 , \427 , \388 );
mxor \mul_6_19_g11475/U$1 ( \429 , \328 , \329 );
mand \mul_6_19_g11436/U$2 ( \430 , \429 , \326 );
mnot \mul_6_19_g11436/U$4 ( \431 , \429 );
mnot \mul_6_19_g11518/U$1 ( \432 , \326 );
mand \mul_6_19_g11436/U$3 ( \433 , \431 , \432 );
mor \mul_6_19_g11436/U$1 ( \434 , \430 , \433 );
mxor \g11855/U$1 ( \435 , \428 , \434 );
mnot \mul_6_19_g11494/U$3 ( \436 , \367 );
mnot \mul_6_19_g11494/U$4 ( \437 , \354 );
mor \mul_6_19_g11494/U$2 ( \438 , \436 , \437 );
mnot \mul_6_19_g11776/U$2 ( \439 , \367 );
mnand \mul_6_19_g11776/U$1 ( \440 , \439 , \352 );
mnand \mul_6_19_g11494/U$1 ( \441 , \438 , \440 );
mand \mul_6_19_g11466/U$2 ( \442 , \441 , \340 );
mnot \mul_6_19_g11466/U$4 ( \443 , \441 );
mnot \fopt11895/U$1 ( \444 , \340 );
mand \mul_6_19_g11466/U$3 ( \445 , \443 , \444 );
mnor \mul_6_19_g11466/U$1 ( \446 , \442 , \445 );
mnand \mul_6_19_g11758/U$1 ( \447 , \80 , \B[4] );
mnand \mul_6_19_g11663/U$1 ( \448 , \88 , \B[2] );
mxor \mul_6_19_g11556/U$4 ( \449 , \447 , \448 );
mnand \mul_6_19_g11664/U$1 ( \450 , \B[9] , \296 );
mand \mul_6_19_g11556/U$3 ( \451 , \449 , \450 );
mand \mul_6_19_g11556/U$5 ( \452 , \447 , \448 );
mor \mul_6_19_g11556/U$2 ( \453 , \451 , \452 );
mxor \mul_6_19_g11759/U$1 ( \454 , \358 , \363 );
mxor \mul_6_19_g11759/U$1_r1 ( \455 , \454 , \360 );
mxor \mul_6_19_g11445/U$4 ( \456 , \453 , \455 );
mand \mul_6_19_g11711/U$1 ( \457 , \119 , \B[3] );
mand \mul_6_19_g11708/U$1 ( \458 , \253 , \B[7] );
mor \mul_6_19_g11787/U$1 ( \459 , \457 , \458 );
mnand \mul_6_19_g11671/U$1 ( \460 , \289 , \B[8] );
mnot \mul_6_19_g11670/U$1 ( \461 , \460 );
mand \mul_6_19_g11537/U$2 ( \462 , \459 , \461 );
mand \mul_6_19_g11576/U$2 ( \463 , \457 , \458 );
mnor \mul_6_19_g11537/U$1 ( \464 , \462 , \463 );
mand \mul_6_19_g11445/U$3 ( \465 , \456 , \464 );
mand \mul_6_19_g11445/U$5 ( \466 , \453 , \455 );
mor \mul_6_19_g11445/U$2 ( \467 , \465 , \466 );
mxor \mul_6_19_g11373/U$4 ( \468 , \446 , \467 );
mxor \g11811/U$1 ( \469 , \342 , \350 );
mxor \g11811/U$1_r1 ( \470 , \469 , \347 );
mnand \mul_6_19_g11626/U$1 ( \471 , \234 , \B[6] );
mnand \mul_6_19_g11643/U$1 ( \472 , \100 , \B[5] );
mxor \mul_6_19_g11507/U$4 ( \473 , \471 , \472 );
mnot \mul_6_19_g11593/U$3 ( \474 , \379 );
mnot \mul_6_19_g11593/U$4 ( \475 , \377 );
mand \mul_6_19_g11593/U$2 ( \476 , \474 , \475 );
mand \mul_6_19_g11593/U$5 ( \477 , \379 , \377 );
mnor \mul_6_19_g11593/U$1 ( \478 , \476 , \477 );
mand \mul_6_19_g11507/U$3 ( \479 , \473 , \478 );
mand \mul_6_19_g11507/U$5 ( \480 , \471 , \472 );
mor \mul_6_19_g11507/U$2 ( \481 , \479 , \480 );
mxor \mul_6_19_g11418/U$4 ( \482 , \470 , \481 );
mand \mul_6_19_g11677/U$1 ( \483 , \88 , \B[0] );
mnand \mul_6_19_g11612/U$1 ( \484 , \379 , \483 );
mnand \mul_6_19_g11683/U$1 ( \485 , \233 , \B[5] );
mnot \mul_6_19_g11582/U$3 ( \486 , \485 );
mnand \mul_6_19_g11700/U$1 ( \487 , \100 , \B[4] );
mnot \mul_6_19_g11582/U$4 ( \488 , \487 );
mor \mul_6_19_g11582/U$2 ( \489 , \486 , \488 );
mand \mul_6_19_g11738/U$1 ( \490 , \119 , \B[2] );
mnand \mul_6_19_g11582/U$1 ( \491 , \489 , \490 );
mnot \mul_6_19_g11599/U$2 ( \492 , \487 );
mnot \mul_6_19_g11682/U$1 ( \493 , \485 );
mnand \mul_6_19_g11599/U$1 ( \494 , \492 , \493 );
mnand \mul_6_19_g11571/U$1 ( \495 , \491 , \494 );
mnot \mul_6_19_g11549/U$1 ( \496 , \495 );
mxor \mul_6_19_g11463/U$4 ( \497 , \484 , \496 );
mnand \mul_6_19_g11752/U$1 ( \498 , \289 , \B[7] );
mnand \mul_6_19_g11673/U$1 ( \499 , \80 , \B[3] );
mnand \mul_6_19_g11616/U$1 ( \500 , \498 , \499 );
mand \mul_6_19_g11648/U$1 ( \501 , \296 , \B[8] );
mand \mul_6_19_g11538/U$2 ( \502 , \500 , \501 );
mnor \mul_6_19_g11614/U$1 ( \503 , \498 , \499 );
mnor \mul_6_19_g11538/U$1 ( \504 , \502 , \503 );
mand \mul_6_19_g11463/U$3 ( \505 , \497 , \504 );
mand \mul_6_19_g11463/U$5 ( \506 , \484 , \496 );
mor \mul_6_19_g11463/U$2 ( \507 , \505 , \506 );
mand \mul_6_19_g11418/U$3 ( \508 , \482 , \507 );
mand \mul_6_19_g11418/U$5 ( \509 , \470 , \481 );
mor \mul_6_19_g11418/U$2 ( \510 , \508 , \509 );
mand \mul_6_19_g11373/U$3 ( \511 , \468 , \510 );
mand \mul_6_19_g11373/U$5 ( \512 , \446 , \467 );
mor \mul_6_19_g11373/U$2 ( \513 , \511 , \512 );
mxnor \mul_6_19_g11334/U$1 ( \514 , \435 , \513 );
mxor \mul_6_19_g11430/U$1 ( \515 , \372 , \374 );
mxor \mul_6_19_g11430/U$1_r1 ( \516 , \515 , \385 );
mxor \mul_6_19_g11487/U$1 ( \517 , \376 , \380 );
mxor \mul_6_19_g11487/U$1_r1 ( \518 , \517 , \382 );
mxor \mul_6_19_g11445/U$1 ( \519 , \453 , \455 );
mxor \mul_6_19_g11445/U$1_r1 ( \520 , \519 , \464 );
mxor \mul_6_19_g11375/U$4 ( \521 , \518 , \520 );
mxor \mul_6_19_g11576/U$1 ( \522 , \457 , \458 );
mand \mul_6_19_g11547/U$2 ( \523 , \522 , \461 );
mnot \mul_6_19_g11547/U$4 ( \524 , \522 );
mand \mul_6_19_g11547/U$3 ( \525 , \524 , \460 );
mnor \mul_6_19_g11547/U$1 ( \526 , \523 , \525 );
mnot \mul_6_19_g11531/U$1 ( \527 , \526 );
mxor \mul_6_19_g11556/U$1 ( \528 , \447 , \448 );
mxor \mul_6_19_g11556/U$1_r1 ( \529 , \528 , \450 );
mnand \mul_6_19_g11502/U$1 ( \530 , \527 , \529 );
mand \mul_6_19_g11696/U$1 ( \531 , \253 , \B[6] );
mand \mul_6_19_g11638/U$1 ( \532 , \88 , \B[1] );
mnot \mul_6_19_g11594/U$3 ( \533 , \532 );
mnand \mul_6_19_g11733/U$1 ( \534 , \140 , \B[0] );
mnot \mul_6_19_g11594/U$4 ( \535 , \534 );
mor \mul_6_19_g11594/U$2 ( \536 , \533 , \535 );
mor \mul_6_19_g11594/U$5 ( \537 , \532 , \534 );
mnand \mul_6_19_g11594/U$1 ( \538 , \536 , \537 );
mxor \mul_6_19_g11486/U$4 ( \539 , \531 , \538 );
mand \mul_6_19_g11741/U$1 ( \540 , \119 , \B[1] );
mand \mul_6_19_g11575/U$2 ( \541 , \483 , \540 );
mand \mul_6_19_g11486/U$3 ( \542 , \539 , \541 );
mand \mul_6_19_g11486/U$5 ( \543 , \531 , \538 );
mor \mul_6_19_g11486/U$2 ( \544 , \542 , \543 );
mand \mul_6_19_g11434/U$2 ( \545 , \530 , \544 );
mnor \mul_6_19_g11501/U$1 ( \546 , \527 , \529 );
mnor \mul_6_19_g11434/U$1 ( \547 , \545 , \546 );
mand \mul_6_19_g11375/U$3 ( \548 , \521 , \547 );
mand \mul_6_19_g11375/U$5 ( \549 , \518 , \520 );
mor \mul_6_19_g11375/U$2 ( \550 , \548 , \549 );
mxor \mul_6_19_g11879/U$4 ( \551 , \516 , \550 );
mxor \mul_6_19_g11373/U$1 ( \552 , \446 , \467 );
mxor \mul_6_19_g11373/U$1_r1 ( \553 , \552 , \510 );
mand \mul_6_19_g11879/U$3 ( \554 , \551 , \553 );
mand \mul_6_19_g11879/U$5 ( \555 , \516 , \550 );
mor \mul_6_19_g11879/U$2 ( \556 , \554 , \555 );
mnand \mul_6_19_g11309/U$1 ( \557 , \514 , \556 );
mnot \mul_6_19_g11339/U$3 ( \558 , \428 );
mnot \mul_6_19_g11427/U$1 ( \559 , \434 );
mnot \mul_6_19_g11339/U$4 ( \560 , \559 );
mor \mul_6_19_g11339/U$2 ( \561 , \558 , \560 );
mnot \mul_6_19_g11372/U$1 ( \562 , \513 );
mnand \mul_6_19_g11339/U$1 ( \563 , \561 , \562 );
mnot \mul_6_19_g11769/U$2 ( \564 , \428 );
mnand \mul_6_19_g11769/U$1 ( \565 , \564 , \434 );
mnand \mul_6_19_g11331/U$1 ( \566 , \563 , \565 );
mnot \mul_6_19_g11765/U$2 ( \567 , \566 );
mxor \mul_6_19_g11841/U$1 ( \568 , \331 , \391 );
mxor \mul_6_19_g11841/U$1_r1 ( \569 , \568 , \334 );
mnand \mul_6_19_g11765/U$1 ( \570 , \567 , \569 );
mnand \mul_6_19_g11294/U$1 ( \571 , \557 , \570 );
mnor \mul_6_19_g11762/U$1 ( \572 , \426 , \571 );
mnot \mul_6_19_g11249/U$3 ( \573 , \572 );
mnand \mul_6_19_g11657/U$1 ( \574 , \119 , \B[0] );
mnot \mul_6_19_g11590/U$3 ( \575 , \574 );
mand \mul_6_19_g11623/U$1 ( \576 , \80 , \B[1] );
mnot \mul_6_19_g11590/U$4 ( \577 , \576 );
mand \mul_6_19_g11590/U$2 ( \578 , \575 , \577 );
mand \mul_6_19_g11590/U$5 ( \579 , \574 , \576 );
mnor \mul_6_19_g11590/U$1 ( \580 , \578 , \579 );
mnand \mul_6_19_g11736/U$1 ( \581 , \289 , \B[4] );
mnand \mul_6_19_g11624/U$1 ( \582 , \234 , \B[2] );
mxor \mul_6_19_g11550/U$4 ( \583 , \581 , \582 );
mnand \mul_6_19_g11743/U$1 ( \584 , \253 , \B[3] );
mand \mul_6_19_g11550/U$3 ( \585 , \583 , \584 );
mand \mul_6_19_g11550/U$5 ( \586 , \581 , \582 );
mor \mul_6_19_g11550/U$2 ( \587 , \585 , \586 );
mxor \mul_6_19_g11465/U$4 ( \588 , \580 , \587 );
mnand \mul_6_19_g11654/U$1 ( \589 , \253 , \B[4] );
mand \mul_6_19_g11760/U$1 ( \590 , \233 , \B[3] );
mxor \g12010/U$1 ( \591 , \589 , \590 );
mnand \mul_6_19_g11732/U$1 ( \592 , \100 , \B[2] );
mxnor \g12010/U$1_r1 ( \593 , \591 , \592 );
mand \mul_6_19_g11465/U$3 ( \594 , \588 , \593 );
mand \mul_6_19_g11465/U$5 ( \595 , \580 , \587 );
mor \mul_6_19_g11465/U$2 ( \596 , \594 , \595 );
mnot \mul_6_19_g11426/U$3 ( \597 , \596 );
mnot \mul_6_19_g11780/U$2 ( \598 , \576 );
mnor \mul_6_19_g11780/U$1 ( \599 , \598 , \574 );
mxor \mul_6_19_g11575/U$1 ( \600 , \483 , \540 );
mxor \mul_6_19_g11478/U$1 ( \601 , \599 , \600 );
mnot \mul_6_19_g11583/U$3 ( \602 , \592 );
mnot \mul_6_19_g11583/U$4 ( \603 , \589 );
mor \mul_6_19_g11583/U$2 ( \604 , \602 , \603 );
mnand \mul_6_19_g11583/U$1 ( \605 , \604 , \590 );
mor \mul_6_19_g11783/U$1 ( \606 , \589 , \592 );
mnand \mul_6_19_g11572/U$1 ( \607 , \605 , \606 );
mxor \mul_6_19_g11478/U$1_r1 ( \608 , \601 , \607 );
mnot \mul_6_19_g11426/U$4 ( \609 , \608 );
mand \mul_6_19_g11426/U$2 ( \610 , \597 , \609 );
mand \mul_6_19_g11426/U$5 ( \611 , \596 , \608 );
mnor \mul_6_19_g11426/U$1 ( \612 , \610 , \611 );
mnand \mul_6_19_g11628/U$1 ( \613 , \80 , \B[2] );
mnand \mul_6_19_g11740/U$1 ( \614 , \253 , \B[5] );
mxor \mul_6_19_g11789/U$1 ( \615 , \613 , \614 );
mnand \mul_6_19_g11666/U$1 ( \616 , \289 , \B[6] );
mxor \mul_6_19_g11789/U$1_r1 ( \617 , \615 , \616 );
mnot \mul_6_19_g11553/U$1 ( \618 , \617 );
mnot \mul_6_19_g11503/U$3 ( \619 , \618 );
mnand \mul_6_19_g11669/U$1 ( \620 , \296 , \B[7] );
mand \g11988/U$1 ( \621 , \100 , \B[3] );
mxor \g11957/U$1 ( \622 , \620 , \621 );
mnand \mul_6_19_g11748/U$1 ( \623 , \234 , \B[4] );
mxnor \g11957/U$1_r1 ( \624 , \622 , \623 );
mnot \mul_6_19_g11503/U$4 ( \625 , \624 );
mor \mul_6_19_g11503/U$2 ( \626 , \619 , \625 );
mnot \mul_6_19_g11551/U$1 ( \627 , \624 );
mnand \mul_6_19_g11504/U$1 ( \628 , \627 , \617 );
mnand \mul_6_19_g11503/U$1 ( \629 , \626 , \628 );
mand \mul_6_19_g11725/U$1 ( \630 , \296 , \B[6] );
mnot \mul_6_19_g11724/U$1 ( \631 , \630 );
mnand \mul_6_19_g11704/U$1 ( \632 , \289 , \B[5] );
mor \mul_6_19_g11540/U$2 ( \633 , \631 , \632 );
mnot \mul_6_19_g11563/U$3 ( \634 , \632 );
mnot \mul_6_19_g11563/U$4 ( \635 , \631 );
mor \mul_6_19_g11563/U$2 ( \636 , \634 , \635 );
mnand \mul_6_19_g11661/U$1 ( \637 , \100 , \B[1] );
mnot \mul_6_19_g11608/U$2 ( \638 , \637 );
mand \mul_6_19_g11713/U$1 ( \639 , \80 , \B[0] );
mnand \mul_6_19_g11608/U$1 ( \640 , \638 , \639 );
mnot \mul_6_19_g11577/U$1 ( \641 , \640 );
mnand \mul_6_19_g11563/U$1 ( \642 , \636 , \641 );
mnand \mul_6_19_g11540/U$1 ( \643 , \633 , \642 );
mnot \mul_6_19_g11511/U$1 ( \644 , \643 );
mand \mul_6_19_g11461/U$2 ( \645 , \629 , \644 );
mnot \mul_6_19_g11461/U$4 ( \646 , \629 );
mand \mul_6_19_g11461/U$3 ( \647 , \646 , \643 );
mnor \mul_6_19_g11461/U$1 ( \648 , \645 , \647 );
mnot \mul_6_19_g11444/U$1 ( \649 , \648 );
mand \mul_6_19_g11405/U$2 ( \650 , \612 , \649 );
mnot \mul_6_19_g11405/U$4 ( \651 , \612 );
mand \mul_6_19_g11405/U$3 ( \652 , \651 , \648 );
mnor \mul_6_19_g11405/U$1 ( \653 , \650 , \652 );
mxor \g11815/U$1 ( \654 , \630 , \632 );
mxnor \g11815/U$1_r1 ( \655 , \654 , \640 );
mnand \mul_6_19_g11726/U$1 ( \656 , \296 , \B[5] );
mnand \mul_6_19_g11698/U$1 ( \657 , \100 , \B[0] );
mnot \mul_6_19_g11613/U$2 ( \658 , \657 );
mand \mul_6_19_g11761/U$1 ( \659 , \233 , \B[1] );
mnand \mul_6_19_g11613/U$1 ( \660 , \658 , \659 );
mxor \mul_6_19_g11489/U$4 ( \661 , \656 , \660 );
mnot \mul_6_19_g11588/U$3 ( \662 , \639 );
mnot \mul_6_19_g11588/U$4 ( \663 , \637 );
mand \mul_6_19_g11588/U$2 ( \664 , \662 , \663 );
mand \mul_6_19_g11588/U$5 ( \665 , \637 , \639 );
mnor \mul_6_19_g11588/U$1 ( \666 , \664 , \665 );
mand \mul_6_19_g11489/U$3 ( \667 , \661 , \666 );
mand \mul_6_19_g11489/U$5 ( \668 , \656 , \660 );
mor \mul_6_19_g11489/U$2 ( \669 , \667 , \668 );
mxor \mul_6_19_g11412/U$4 ( \670 , \655 , \669 );
mxor \mul_6_19_g11465/U$1 ( \671 , \580 , \587 );
mxor \mul_6_19_g11465/U$1_r1 ( \672 , \671 , \593 );
mand \mul_6_19_g11412/U$3 ( \673 , \670 , \672 );
mand \mul_6_19_g11412/U$5 ( \674 , \655 , \669 );
mor \mul_6_19_g11412/U$2 ( \675 , \673 , \674 );
mnand \mul_6_19_g11381/U$1 ( \676 , \653 , \675 );
mnot \mul_6_19_g11320/U$3 ( \677 , \676 );
mxor \mul_6_19_g11412/U$1 ( \678 , \655 , \669 );
mxor \mul_6_19_g11412/U$1_r1 ( \679 , \678 , \672 );
mnand \mul_6_19_g11642/U$1 ( \680 , \296 , \B[4] );
mnand \mul_6_19_g11678/U$1 ( \681 , \253 , \B[2] );
mxor \mul_6_19_g11557/U$4 ( \682 , \680 , \681 );
mnand \mul_6_19_g11639/U$1 ( \683 , \289 , \B[3] );
mand \mul_6_19_g11557/U$3 ( \684 , \682 , \683 );
mand \mul_6_19_g11557/U$5 ( \685 , \680 , \681 );
mor \mul_6_19_g11557/U$2 ( \686 , \684 , \685 );
mxor \mul_6_19_g11550/U$1 ( \687 , \581 , \582 );
mxor \mul_6_19_g11550/U$1_r1 ( \688 , \687 , \584 );
mxor \mul_6_19_g11448/U$4 ( \689 , \686 , \688 );
mxor \mul_6_19_g11489/U$1 ( \690 , \656 , \660 );
mxor \mul_6_19_g11489/U$1_r1 ( \691 , \690 , \666 );
mand \mul_6_19_g11448/U$3 ( \692 , \689 , \691 );
mand \mul_6_19_g11448/U$5 ( \693 , \686 , \688 );
mor \mul_6_19_g11448/U$2 ( \694 , \692 , \693 );
mnand \mul_6_19_g11397/U$1 ( \695 , \679 , \694 );
mnot \mul_6_19_g11350/U$3 ( \696 , \695 );
mxor \mul_6_19_g11448/U$1 ( \697 , \686 , \688 );
mxor \mul_6_19_g11448/U$1_r1 ( \698 , \697 , \691 );
mnand \mul_6_19_g11652/U$1 ( \699 , \234 , \B[0] );
mnot \mul_6_19_g11782/U$2 ( \700 , \699 );
mand \mul_6_19_g11684/U$1 ( \701 , \253 , \B[1] );
mnand \mul_6_19_g11782/U$1 ( \702 , \700 , \701 );
mnot \mul_6_19_g11591/U$3 ( \703 , \659 );
mnot \mul_6_19_g11591/U$4 ( \704 , \657 );
mand \mul_6_19_g11591/U$2 ( \705 , \703 , \704 );
mand \mul_6_19_g11591/U$5 ( \706 , \659 , \657 );
mnor \mul_6_19_g11591/U$1 ( \707 , \705 , \706 );
mxor \mul_6_19_g11481/U$4 ( \708 , \702 , \707 );
mxor \mul_6_19_g11557/U$1 ( \709 , \680 , \681 );
mxor \mul_6_19_g11557/U$1_r1 ( \710 , \709 , \683 );
mand \mul_6_19_g11481/U$3 ( \711 , \708 , \710 );
mand \mul_6_19_g11481/U$5 ( \712 , \702 , \707 );
mor \mul_6_19_g11481/U$2 ( \713 , \711 , \712 );
mnand \mul_6_19_g11423/U$1 ( \714 , \698 , \713 );
mnot \mul_6_19_g11385/U$3 ( \715 , \714 );
mxor \mul_6_19_g11481/U$1 ( \716 , \702 , \707 );
mxor \mul_6_19_g11481/U$1_r1 ( \717 , \716 , \710 );
mnot \mul_6_19_g11592/U$3 ( \718 , \701 );
mnot \mul_6_19_g11592/U$4 ( \719 , \699 );
mand \mul_6_19_g11592/U$2 ( \720 , \718 , \719 );
mand \mul_6_19_g11592/U$5 ( \721 , \699 , \701 );
mnor \mul_6_19_g11592/U$1 ( \722 , \720 , \721 );
mnot \g11865/U$2 ( \723 , \722 );
mand \mul_6_19_g11620/U$1 ( \724 , \296 , \B[3] );
mnot \g11866/U$2 ( \725 , \724 );
mnand \mul_6_19_g11705/U$1 ( \726 , \289 , \B[2] );
mnand \g11866/U$1 ( \727 , \725 , \726 );
mnand \g11865/U$1 ( \728 , \723 , \727 );
mnot \mul_6_19_g11607/U$2 ( \729 , \726 );
mnand \mul_6_19_g11607/U$1 ( \730 , \729 , \724 );
mand \mul_6_19_g11539/U$1 ( \731 , \728 , \730 );
mor \mul_6_19_g11773/U$1 ( \732 , \717 , \731 );
mand \mul_6_19_g11729/U$1 ( \733 , \253 , \B[0] );
mand \mul_6_19_g11646/U$1 ( \734 , \296 , \B[2] );
mand \mul_6_19_g11574/U$2 ( \735 , \733 , \734 );
mnot \mul_6_19_g11779/U$2 ( \736 , \735 );
mnot \mul_6_19_g11546/U$3 ( \737 , \722 );
mnot \mul_6_19_g11597/U$3 ( \738 , \726 );
mnot \mul_6_19_g11597/U$4 ( \739 , \724 );
mor \mul_6_19_g11597/U$2 ( \740 , \738 , \739 );
mor \mul_6_19_g11597/U$5 ( \741 , \724 , \726 );
mnand \mul_6_19_g11597/U$1 ( \742 , \740 , \741 );
mnot \mul_6_19_g11546/U$4 ( \743 , \742 );
mand \mul_6_19_g11546/U$2 ( \744 , \737 , \743 );
mand \mul_6_19_g11546/U$5 ( \745 , \742 , \722 );
mnor \mul_6_19_g11546/U$1 ( \746 , \744 , \745 );
mnand \mul_6_19_g11779/U$1 ( \747 , \736 , \746 );
mnot \g11955/U$3 ( \748 , \747 );
mnand \mul_6_19_g11691/U$1 ( \749 , \289 , \B[1] );
mnot \mul_6_19_g11690/U$1 ( \750 , \749 );
mnand \mul_6_19_g11645/U$1 ( \751 , \296 , \B[0] );
mnor \mul_6_19_g11615/U$1 ( \752 , \749 , \751 );
mxor \mul_6_19_g11484/U$4 ( \753 , \750 , \752 );
mxor \mul_6_19_g11574/U$1 ( \754 , \733 , \734 );
mand \mul_6_19_g11484/U$3 ( \755 , \753 , \754 );
mand \mul_6_19_g11484/U$5 ( \756 , \750 , \752 );
mor \mul_6_19_g11484/U$2 ( \757 , \755 , \756 );
mnot \g11955/U$4 ( \758 , \757 );
mor \g11955/U$2 ( \759 , \748 , \758 );
mnot \mul_6_19_g11777/U$2 ( \760 , \746 );
mnand \mul_6_19_g11777/U$1 ( \761 , \760 , \735 );
mnand \g11955/U$1 ( \762 , \759 , \761 );
mnand \mul_6_19_g11453/U$1 ( \763 , \717 , \731 );
mnand \mul_6_19_g11424/U$1 ( \764 , \762 , \763 );
mnand \mul_6_19_g11416/U$1 ( \765 , \732 , \764 );
mnot \mul_6_19_g11385/U$4 ( \766 , \765 );
mor \mul_6_19_g11385/U$2 ( \767 , \715 , \766 );
mor \mul_6_19_g11772/U$1 ( \768 , \698 , \713 );
mnand \mul_6_19_g11385/U$1 ( \769 , \767 , \768 );
mnot \mul_6_19_g11350/U$4 ( \770 , \769 );
mor \mul_6_19_g11350/U$2 ( \771 , \696 , \770 );
mnot \mul_6_19_g11410/U$1 ( \772 , \679 );
mnot \mul_6_19_g11447/U$1 ( \773 , \694 );
mnand \mul_6_19_g11396/U$1 ( \774 , \772 , \773 );
mnand \mul_6_19_g11350/U$1 ( \775 , \771 , \774 );
mnot \mul_6_19_g11320/U$4 ( \776 , \775 );
mor \mul_6_19_g11320/U$2 ( \777 , \677 , \776 );
mnot \mul_6_19_g11400/U$1 ( \778 , \653 );
mnot \mul_6_19_g11411/U$1 ( \779 , \675 );
mnand \mul_6_19_g11380/U$1 ( \780 , \778 , \779 );
mnand \mul_6_19_g11320/U$1 ( \781 , \777 , \780 );
mnot \mul_6_19_g11470/U$3 ( \782 , \617 );
mnot \mul_6_19_g11470/U$4 ( \783 , \624 );
mor \mul_6_19_g11470/U$2 ( \784 , \782 , \783 );
mnand \mul_6_19_g11470/U$1 ( \785 , \784 , \643 );
mnand \mul_6_19_g11505/U$1 ( \786 , \627 , \618 );
mnand \mul_6_19_g11458/U$1 ( \787 , \785 , \786 );
mnot \mul_6_19_g11581/U$3 ( \788 , \623 );
mnot \mul_6_19_g11581/U$4 ( \789 , \620 );
mor \mul_6_19_g11581/U$2 ( \790 , \788 , \789 );
mnand \mul_6_19_g11581/U$1 ( \791 , \790 , \621 );
mor \mul_6_19_g11786/U$1 ( \792 , \623 , \620 );
mnand \mul_6_19_g11569/U$1 ( \793 , \791 , \792 );
mnot \mul_6_19_g11580/U$3 ( \794 , \614 );
mnot \mul_6_19_g11580/U$4 ( \795 , \616 );
mor \mul_6_19_g11580/U$2 ( \796 , \794 , \795 );
mnot \mul_6_19_g11627/U$1 ( \797 , \613 );
mnand \mul_6_19_g11580/U$1 ( \798 , \796 , \797 );
mor \mul_6_19_g11785/U$1 ( \799 , \614 , \616 );
mnand \mul_6_19_g11570/U$1 ( \800 , \798 , \799 );
mxor \mul_6_19_g11488/U$1 ( \801 , \793 , \800 );
mxor \g12023/U$1 ( \802 , \490 , \487 );
mnot \g12023/U$2 ( \803 , \485 );
mxor \g12023/U$1_r1 ( \804 , \802 , \803 );
mnot \mul_6_19_g11548/U$1 ( \805 , \804 );
mand \mul_6_19_g11462/U$2 ( \806 , \801 , \805 );
mnot \mul_6_19_g11462/U$4 ( \807 , \801 );
mand \mul_6_19_g11462/U$3 ( \808 , \807 , \804 );
mnor \mul_6_19_g11462/U$1 ( \809 , \806 , \808 );
mxor \mul_6_19_g11379/U$1 ( \810 , \787 , \809 );
mxor \mul_6_19_g11541/U$1 ( \811 , \499 , \498 );
mxor \mul_6_19_g11541/U$1_r1 ( \812 , \811 , \501 );
mxor \mul_6_19_g11486/U$1 ( \813 , \531 , \538 );
mxor \mul_6_19_g11486/U$1_r1 ( \814 , \813 , \541 );
mxor \mul_6_19_g11409/U$1 ( \815 , \812 , \814 );
mxor \mul_6_19_g11478/U$4 ( \816 , \599 , \600 );
mand \mul_6_19_g11478/U$3 ( \817 , \816 , \607 );
mand \mul_6_19_g11478/U$5 ( \818 , \599 , \600 );
mor \mul_6_19_g11478/U$2 ( \819 , \817 , \818 );
mxor \mul_6_19_g11409/U$1_r1 ( \820 , \815 , \819 );
mxor \mul_6_19_g11379/U$1_r1 ( \821 , \810 , \820 );
mnot \mul_6_19_g11377/U$1 ( \822 , \821 );
mnot \g11953/U$3 ( \823 , \608 );
mnot \g11953/U$4 ( \824 , \649 );
mor \g11953/U$2 ( \825 , \823 , \824 );
mnot \mul_6_19_g11954/U$1 ( \826 , \608 );
mnot \mul_6_19_g11414/U$3 ( \827 , \826 );
mnot \mul_6_19_g11414/U$4 ( \828 , \648 );
mor \mul_6_19_g11414/U$2 ( \829 , \827 , \828 );
mnot \mul_6_19_g11464/U$1 ( \830 , \596 );
mnand \mul_6_19_g11414/U$1 ( \831 , \829 , \830 );
mnand \g11953/U$1 ( \832 , \825 , \831 );
mnot \mul_6_19_g11401/U$1 ( \833 , \832 );
mnand \mul_6_19_g11361/U$1 ( \834 , \822 , \833 );
mnand \mul_6_19_g11285/U$1 ( \835 , \781 , \834 );
mand \g12008/U$2 ( \836 , \529 , \526 );
mnot \g12008/U$4 ( \837 , \529 );
mand \g12008/U$3 ( \838 , \837 , \527 );
mor \g12008/U$1 ( \839 , \836 , \838 );
mxor \mul_6_19_g11774/U$1 ( \840 , \839 , \544 );
mxor \mul_6_19_g11409/U$4 ( \841 , \812 , \814 );
mand \mul_6_19_g11409/U$3 ( \842 , \841 , \819 );
mand \mul_6_19_g11409/U$5 ( \843 , \812 , \814 );
mor \mul_6_19_g11409/U$2 ( \844 , \842 , \843 );
mxor \mul_6_19_g11376/U$1 ( \845 , \840 , \844 );
mxor \mul_6_19_g11507/U$1 ( \846 , \471 , \472 );
mxor \mul_6_19_g11507/U$1_r1 ( \847 , \846 , \478 );
mxor \mul_6_19_g11463/U$1 ( \848 , \484 , \496 );
mxor \mul_6_19_g11463/U$1_r1 ( \849 , \848 , \504 );
mxor \mul_6_19_g11391/U$1 ( \850 , \847 , \849 );
mor \mul_6_19_g11778/U$1 ( \851 , \793 , \800 );
mand \mul_6_19_g11457/U$2 ( \852 , \851 , \805 );
mand \mul_6_19_g11488/U$2 ( \853 , \793 , \800 );
mnor \mul_6_19_g11457/U$1 ( \854 , \852 , \853 );
mxor \mul_6_19_g11391/U$1_r1 ( \855 , \850 , \854 );
mnot \mul_6_19_g11388/U$1 ( \856 , \855 );
mand \mul_6_19_g11351/U$2 ( \857 , \845 , \856 );
mnot \mul_6_19_g11351/U$4 ( \858 , \845 );
mand \mul_6_19_g11351/U$3 ( \859 , \858 , \855 );
mnor \mul_6_19_g11351/U$1 ( \860 , \857 , \859 );
mxor \mul_6_19_g11379/U$4 ( \861 , \787 , \809 );
mand \mul_6_19_g11379/U$3 ( \862 , \861 , \820 );
mand \mul_6_19_g11379/U$5 ( \863 , \787 , \809 );
mor \mul_6_19_g11379/U$2 ( \864 , \862 , \863 );
mnand \mul_6_19_g11327/U$1 ( \865 , \860 , \864 );
mnand \mul_6_19_g11360/U$1 ( \866 , \821 , \832 );
mand \mul_6_19_g11314/U$1 ( \867 , \865 , \866 );
mnand \mul_6_19_g11281/U$1 ( \868 , \835 , \867 );
mnot \mul_6_19_g11265/U$3 ( \869 , \868 );
mxor \mul_6_19_g11418/U$1 ( \870 , \470 , \481 );
mxor \mul_6_19_g11418/U$1_r1 ( \871 , \870 , \507 );
mnot \mul_6_19_g11363/U$3 ( \872 , \871 );
mxor \mul_6_19_g11391/U$4 ( \873 , \847 , \849 );
mand \mul_6_19_g11391/U$3 ( \874 , \873 , \854 );
mand \mul_6_19_g11391/U$5 ( \875 , \847 , \849 );
mor \mul_6_19_g11391/U$2 ( \876 , \874 , \875 );
mnot \mul_6_19_g11390/U$1 ( \877 , \876 );
mnot \mul_6_19_g11363/U$4 ( \878 , \877 );
mor \mul_6_19_g11363/U$2 ( \879 , \872 , \878 );
mnot \mul_6_19_g11365/U$2 ( \880 , \871 );
mnand \mul_6_19_g11365/U$1 ( \881 , \880 , \876 );
mnand \mul_6_19_g11363/U$1 ( \882 , \879 , \881 );
mxor \mul_6_19_g11375/U$1 ( \883 , \518 , \520 );
mxor \mul_6_19_g11375/U$1_r1 ( \884 , \883 , \547 );
mxor \g11859/U$1 ( \885 , \882 , \884 );
mor \mul_6_19_g11770/U$1 ( \886 , \844 , \840 );
mand \mul_6_19_g11349/U$2 ( \887 , \856 , \886 );
mand \mul_6_19_g11376/U$2 ( \888 , \840 , \844 );
mnor \mul_6_19_g11349/U$1 ( \889 , \887 , \888 );
mnand \mul_6_19_g11317/U$1 ( \890 , \885 , \889 );
mnot \mul_6_19_g11328/U$2 ( \891 , \860 );
mnot \mul_6_19_g11378/U$1 ( \892 , \864 );
mnand \mul_6_19_g11328/U$1 ( \893 , \891 , \892 );
mnand \mul_6_19_g11305/U$1 ( \894 , \890 , \893 );
mxor \g11878/U$1 ( \895 , \516 , \550 );
mxnor \g11878/U$1_r1 ( \896 , \895 , \553 );
mnot \mul_6_19_g11348/U$3 ( \897 , \871 );
mnot \mul_6_19_g11348/U$4 ( \898 , \884 );
mor \mul_6_19_g11348/U$2 ( \899 , \897 , \898 );
mnot \mul_6_19_g11389/U$1 ( \900 , \876 );
mnand \mul_6_19_g11348/U$1 ( \901 , \899 , \900 );
mnot \mul_6_19_g11362/U$2 ( \902 , \871 );
mnot \mul_6_19_g11860/U$1 ( \903 , \884 );
mnand \mul_6_19_g11362/U$1 ( \904 , \902 , \903 );
mnand \mul_6_19_g11341/U$1 ( \905 , \901 , \904 );
mnor \mul_6_19_g11297/U$1 ( \906 , \896 , \905 );
mnor \mul_6_19_g11295/U$1 ( \907 , \894 , \906 );
mnot \mul_6_19_g11265/U$4 ( \908 , \907 );
mor \mul_6_19_g11265/U$2 ( \909 , \869 , \908 );
mxor \mul_6_19_g11879/U$1 ( \910 , \516 , \550 );
mxor \mul_6_19_g11879/U$1_r1 ( \911 , \910 , \553 );
mnot \mul_6_19_g11335/U$1 ( \912 , \905 );
mnand \mul_6_19_g11298/U$1 ( \913 , \911 , \912 );
mnor \mul_6_19_g11313/U$1 ( \914 , \885 , \889 );
mand \mul_6_19_g11280/U$2 ( \915 , \913 , \914 );
mnor \mul_6_19_g11310/U$1 ( \916 , \911 , \912 );
mnor \mul_6_19_g11280/U$1 ( \917 , \915 , \916 );
mnand \mul_6_19_g11265/U$1 ( \918 , \909 , \917 );
mnot \mul_6_19_g11249/U$4 ( \919 , \918 );
mor \mul_6_19_g11249/U$2 ( \920 , \573 , \919 );
mnot \mul_6_19_g11279/U$3 ( \921 , \570 );
mnor \mul_6_19_g11304/U$1 ( \922 , \514 , \556 );
mnot \mul_6_19_g11279/U$4 ( \923 , \922 );
mor \mul_6_19_g11279/U$2 ( \924 , \921 , \923 );
mnot \mul_6_19_g11763/U$2 ( \925 , \569 );
mnand \mul_6_19_g11763/U$1 ( \926 , \925 , \566 );
mnand \mul_6_19_g11279/U$1 ( \927 , \924 , \926 );
mnand \mul_6_19_g11268/U$1 ( \928 , \927 , \425 );
mnot \mul_6_19_g11767/U$2 ( \929 , \423 );
mnand \mul_6_19_g11306/U$1 ( \930 , \395 , \397 );
mnor \mul_6_19_g11286/U$1 ( \931 , \930 , \271 );
mnor \mul_6_19_g11275/U$1 ( \932 , \931 , \275 );
mnor \mul_6_19_g11767/U$1 ( \933 , \929 , \932 );
mnor \mul_6_19_g11359/U$1 ( \934 , \420 , \422 );
mor \mul_6_19_g11261/U$2 ( \935 , \933 , \934 );
mnand \mul_6_19_g11261/U$1 ( \936 , \935 , \416 );
mor \mul_6_19_g11398/U$1 ( \937 , \413 , \415 );
mand \mul_6_19_g11255/U$1 ( \938 , \928 , \936 , \937 );
mnand \mul_6_19_g11249/U$1 ( \939 , \920 , \938 );
mnot \mul_6_19_g11245/U$4 ( \940 , \939 );
mor \mul_6_19_g11245/U$2 ( \941 , \312 , \940 );
mor \mul_6_19_g11451/U$1 ( \942 , \309 , \310 );
mnand \mul_6_19_g11245/U$1 ( \943 , \941 , \942 );
mnand \mul_6_19_g11431/U$1 ( \944 , \311 , \942 );
mnot \mul_6_19_g11246/U$3 ( \945 , \944 );
mnot \mul_6_19_g11246/U$4 ( \946 , \939 );
mor \mul_6_19_g11246/U$2 ( \947 , \945 , \946 );
mor \mul_6_19_g11246/U$5 ( \948 , \944 , \939 );
mnand \mul_6_19_g11246/U$1 ( \949 , \947 , \948 );
mnot \mul_6_19_g11250/U$3 ( \950 , \423 );
mnor \mul_6_19_g11272/U$1 ( \951 , \571 , \399 );
mnot \mul_6_19_g11258/U$3 ( \952 , \951 );
mnot \mul_6_19_g11258/U$4 ( \953 , \918 );
mor \mul_6_19_g11258/U$2 ( \954 , \952 , \953 );
mand \g11857/U$1 ( \955 , \398 , \272 );
mand \mul_6_19_g11264/U$2 ( \956 , \927 , \955 );
mnot \mul_6_19_g11274/U$1 ( \957 , \932 );
mnor \mul_6_19_g11264/U$1 ( \958 , \956 , \957 );
mnand \mul_6_19_g11258/U$1 ( \959 , \954 , \958 );
mnot \mul_6_19_g11250/U$4 ( \960 , \959 );
mor \mul_6_19_g11250/U$2 ( \961 , \950 , \960 );
mnot \mul_6_19_g11358/U$1 ( \962 , \934 );
mnand \mul_6_19_g11250/U$1 ( \963 , \961 , \962 );
mnand \mul_6_19_g11384/U$1 ( \964 , \416 , \937 );
mnot \mul_6_19_g11383/U$1 ( \965 , \964 );
mand \mul_6_19_g11247/U$2 ( \966 , \963 , \965 );
mnot \mul_6_19_g11247/U$4 ( \967 , \963 );
mand \mul_6_19_g11247/U$3 ( \968 , \967 , \964 );
mnor \mul_6_19_g11247/U$1 ( \969 , \966 , \968 );
mbuf \fopt11922/U$1 ( \970 , \398 );
mnot \mul_6_19_g11251/U$3 ( \971 , \970 );
mnot \mul_6_19_g11293/U$1 ( \972 , \571 );
mnot \mul_6_19_g11257/U$3 ( \973 , \972 );
mnot \mul_6_19_g11257/U$4 ( \974 , \918 );
mor \mul_6_19_g11257/U$2 ( \975 , \973 , \974 );
mnot \fopt/U$1 ( \976 , \927 );
mnand \mul_6_19_g11257/U$1 ( \977 , \975 , \976 );
mnot \mul_6_19_g11251/U$4 ( \978 , \977 );
mor \mul_6_19_g11251/U$2 ( \979 , \971 , \978 );
mbuf \fopt11892/U$1 ( \980 , \930 );
mnand \mul_6_19_g11251/U$1 ( \981 , \979 , \980 );
mand \mul_6_19_g11248/U$2 ( \982 , \981 , \276 );
mnot \mul_6_19_g11248/U$4 ( \983 , \981 );
mand \mul_6_19_g11248/U$3 ( \984 , \983 , \282 );
mnor \mul_6_19_g11248/U$1 ( \985 , \982 , \984 );
mbuf \fopt11921/U$1 ( \986 , \557 );
mnot \mul_6_19_g11259/U$3 ( \987 , \986 );
mnot \mul_6_19_g11259/U$4 ( \988 , \918 );
mor \mul_6_19_g11259/U$2 ( \989 , \987 , \988 );
mnot \mul_6_19_g11303/U$1 ( \990 , \922 );
mnand \mul_6_19_g11259/U$1 ( \991 , \989 , \990 );
mnand \mul_6_19_g11289/U$1 ( \992 , \570 , \926 );
mnot \mul_6_19_g11288/U$1 ( \993 , \992 );
mand \mul_6_19_g11254/U$2 ( \994 , \991 , \993 );
mnot \mul_6_19_g11254/U$4 ( \995 , \991 );
mand \mul_6_19_g11254/U$3 ( \996 , \995 , \992 );
mnor \mul_6_19_g11254/U$1 ( \997 , \994 , \996 );
mnand \mul_6_19_g11270/U$1 ( \998 , \868 , \893 );
mnot \mul_6_19_g11269/U$1 ( \999 , \998 );
mbuf \mul_6_19_g11316/U$1 ( \1000 , \890 );
mand \mul_6_19_g11262/U$2 ( \1001 , \999 , \1000 );
mbuf \fopt11900/U$1 ( \1002 , \914 );
mnor \mul_6_19_g11262/U$1 ( \1003 , \1001 , \1002 );
mnot \mul_6_19_g11292/U$2 ( \1004 , \916 );
mnand \mul_6_19_g11292/U$1 ( \1005 , \1004 , \913 );
mand \mul_6_19_g11256/U$2 ( \1006 , \1003 , \1005 );
mnot \mul_6_19_g11256/U$4 ( \1007 , \1003 );
mnot \mul_6_19_g11291/U$1 ( \1008 , \1005 );
mand \mul_6_19_g11256/U$3 ( \1009 , \1007 , \1008 );
mnor \mul_6_19_g11256/U$1 ( \1010 , \1006 , \1009 );
mnot \fopt11899/U$1 ( \1011 , \1002 );
mnand \mul_6_19_g11308/U$1 ( \1012 , \1011 , \1000 );
mand \mul_6_19_g11263/U$2 ( \1013 , \998 , \1012 );
mnot \mul_6_19_g11263/U$4 ( \1014 , \998 );
mnot \mul_6_19_g11307/U$1 ( \1015 , \1012 );
mand \mul_6_19_g11263/U$3 ( \1016 , \1014 , \1015 );
mnor \mul_6_19_g11263/U$1 ( \1017 , \1013 , \1016 );
mnand \mul_6_19_g11273/U$1 ( \1018 , \835 , \866 );
mnand \mul_6_19_g11319/U$1 ( \1019 , \893 , \865 );
mnot \mul_6_19_g11318/U$1 ( \1020 , \1019 );
mand \mul_6_19_g11266/U$2 ( \1021 , \1018 , \1020 );
mnot \mul_6_19_g11266/U$4 ( \1022 , \1018 );
mand \mul_6_19_g11266/U$3 ( \1023 , \1022 , \1019 );
mnor \mul_6_19_g11266/U$1 ( \1024 , \1021 , \1023 );
mnand \mul_6_19_g11346/U$1 ( \1025 , \834 , \866 );
mnot \mul_6_19_g11345/U$1 ( \1026 , \1025 );
mand \mul_6_19_g11282/U$2 ( \1027 , \781 , \1026 );
mnot \mul_6_19_g11282/U$4 ( \1028 , \781 );
mand \mul_6_19_g11282/U$3 ( \1029 , \1028 , \1025 );
mnor \mul_6_19_g11282/U$1 ( \1030 , \1027 , \1029 );
mnand \mul_6_19_g11287/U$1 ( \1031 , \970 , \980 );
mnand \mul_6_19_g11290/U$1 ( \1032 , \990 , \986 );
mnand \mul_6_19_g11368/U$1 ( \1033 , \780 , \676 );
mnot \mul_6_19_g11321/U$3 ( \1034 , \1033 );
mbuf \mul_6_19_g11342/U$1 ( \1035 , \775 );
mnot \mul_6_19_g11321/U$4 ( \1036 , \1035 );
mor \mul_6_19_g11321/U$2 ( \1037 , \1034 , \1036 );
mor \mul_6_19_g11321/U$5 ( \1038 , \1035 , \1033 );
mnand \mul_6_19_g11321/U$1 ( \1039 , \1037 , \1038 );
mnand \mul_6_19_g11347/U$1 ( \1040 , \423 , \962 );
mbuf \mul_6_19_g11369/U$1 ( \1041 , \769 );
mnot \mul_6_19_g11352/U$3 ( \1042 , \1041 );
mnand \mul_6_19_g11382/U$1 ( \1043 , \774 , \695 );
mnot \mul_6_19_g11352/U$4 ( \1044 , \1043 );
mor \mul_6_19_g11352/U$2 ( \1045 , \1042 , \1044 );
mor \mul_6_19_g11352/U$5 ( \1046 , \1041 , \1043 );
mnand \mul_6_19_g11352/U$1 ( \1047 , \1045 , \1046 );
mand \mul_6_19_g11771/U$1 ( \1048 , \768 , \714 );
mand \mul_6_19_g11386/U$2 ( \1049 , \1048 , \765 );
mnot \mul_6_19_g11386/U$4 ( \1050 , \1048 );
mnot \mul_6_19_g11406/U$1 ( \1051 , \765 );
mand \mul_6_19_g11386/U$3 ( \1052 , \1050 , \1051 );
mnor \mul_6_19_g11386/U$1 ( \1053 , \1049 , \1052 );
mnand \mul_6_19_g11432/U$1 ( \1054 , \732 , \763 );
mnot \mul_6_19_g11437/U$1 ( \1055 , \762 );
mand \mul_6_19_g11417/U$2 ( \1056 , \1054 , \1055 );
mnot \mul_6_19_g11417/U$4 ( \1057 , \1054 );
mand \mul_6_19_g11417/U$3 ( \1058 , \1057 , \762 );
mnor \mul_6_19_g11417/U$1 ( \1059 , \1056 , \1058 );
mnand \mul_6_19_g11483/U$1 ( \1060 , \761 , \747 );
mnot \mul_6_19_g11460/U$3 ( \1061 , \1060 );
mnot \mul_6_19_g11460/U$4 ( \1062 , \757 );
mor \mul_6_19_g11460/U$2 ( \1063 , \1061 , \1062 );
mor \mul_6_19_g11460/U$5 ( \1064 , \757 , \1060 );
mnand \mul_6_19_g11460/U$1 ( \1065 , \1063 , \1064 );
mxor \mul_6_19_g11484/U$1 ( \1066 , \750 , \752 );
mxor \mul_6_19_g11484/U$1_r1 ( \1067 , \1066 , \754 );
mand \mul_6_19_g11618/U$2 ( \1068 , \289 , \B[0] );
mand \mul_6_19_g11618/U$3 ( \1069 , \296 , \B[1] );
mnor \mul_6_19_g11618/U$1 ( \1070 , \1068 , \1069 );
mnor \mul_6_19_g11579/U$1 ( \1071 , \752 , \1070 );
mnot \mul_6_19_g11644/U$1 ( \1072 , \751 );
mxnor \g2/U$1 ( \1073 , \959 , \1040 );
mxnor \g11791/U$1 ( \1074 , \977 , \1031 );
mxnor \g11792/U$1 ( \1075 , \1032 , \918 );
endmodule


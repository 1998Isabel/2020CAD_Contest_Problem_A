//
// Conformal-LEC Version 19.20-d218 (25-Feb-2020)
//
module top(C, D, O);
input C,D;
output O;


or \g11877/U$2 ( O, C, D );
endmodule


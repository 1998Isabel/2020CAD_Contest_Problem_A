//
// Conformal-LEC Version 19.20-d255 (16-Apr-2020)
//
module top(\a[15] ,\a[14] ,\a[13] ,\a[12] ,\a[11] ,\a[10] ,\a[9] ,\a[8] ,\a[7] ,
        \a[6] ,\a[5] ,\a[4] ,\a[3] ,\a[2] ,\a[1] ,\a[0] ,\b[15] ,\b[14] ,\b[13] ,
        \b[12] ,\b[11] ,\b[10] ,\b[9] ,\b[8] ,\b[7] ,\b[6] ,\b[5] ,\b[4] ,\b[3] ,
        \b[2] ,\b[1] ,\b[0] ,\c[15] ,\c[14] ,\c[13] ,\c[12] ,\c[11] ,\c[10] ,\c[9] ,
        \c[8] ,\c[7] ,\c[6] ,\c[5] ,\c[4] ,\c[3] ,\c[2] ,\c[1] ,\c[0] ,\d[15] ,
        \d[14] ,\d[13] ,\d[12] ,\d[11] ,\d[10] ,\d[9] ,\d[8] ,\d[7] ,\d[6] ,\d[5] ,
        \d[4] ,\d[3] ,\d[2] ,\d[1] ,\d[0] ,\o[31] ,\o[30] ,\o[29] ,\o[28] ,\o[27] ,
        \o[26] ,\o[25] ,\o[24] ,\o[23] ,\o[22] ,\o[21] ,\o[20] ,\o[19] ,\o[18] ,\o[17] ,
        \o[16] ,\o[15] ,\o[14] ,\o[13] ,\o[12] ,\o[11] ,\o[10] ,\o[9] ,\o[8] ,\o[7] ,
        \o[6] ,\o[5] ,\o[4] ,\o[3] ,\o[2] ,\o[1] ,\o[0] );
input [1:0] \a[15] ,\a[14] ,\a[13] ,\a[12] ,\a[11] ,\a[10] ,\a[9] ,\a[8] ,\a[7] ,        \a[6] ,\a[5] ,\a[4] ,\a[3] ,\a[2] ,\a[1] ,\a[0] ,\b[15] ,\b[14] ,\b[13] ,        \b[12] ,\b[11] ,\b[10] ,\b[9] ,\b[8] ,\b[7] ,\b[6] ,\b[5] ,\b[4] ,\b[3] ,        \b[2] ,\b[1] ,\b[0] ,\c[15] ,\c[14] ,\c[13] ,\c[12] ,\c[11] ,\c[10] ,\c[9] ,        \c[8] ,\c[7] ,\c[6] ,\c[5] ,\c[4] ,\c[3] ,\c[2] ,\c[1] ,\c[0] ,\d[15] ,        \d[14] ,\d[13] ,\d[12] ,\d[11] ,\d[10] ,\d[9] ,\d[8] ,\d[7] ,\d[6] ,\d[5] ,        \d[4] ,\d[3] ,\d[2] ,\d[1] ,\d[0] ;
output [1:0] \o[31] ,\o[30] ,\o[29] ,\o[28] ,\o[27] ,\o[26] ,\o[25] ,\o[24] ,\o[23] ,        \o[22] ,\o[21] ,\o[20] ,\o[19] ,\o[18] ,\o[17] ,\o[16] ,\o[15] ,\o[14] ,\o[13] ,        \o[12] ,\o[11] ,\o[10] ,\o[9] ,\o[8] ,\o[7] ,\o[6] ,\o[5] ,\o[4] ,\o[3] ,        \o[2] ,\o[1] ,\o[0] ;

wire [1:0] \97_n22[15] , \98_n22[14] , \99_n22[13] , \100_n22[12] , \101_n22[11] , \102_n22[10] , \103_n22[9] , \104_n22[8] , \105_n22[7] ,         \106_n22[6] , \107_n22[5] , \108_n22[4] , \109_n22[3] , \110_n22[2] , \111_n22[1] , \112_n22[0] , \113_ZERO , \114_ZERO , \115 ,         \116 , \117 , \118 , \119 , \120 , \121 , \122 , \123 , \124 , \125 ,         \126 , \127 , \128 , \129 , \130 , \131 , \132 , \133 , \134 , \135 ,         \136 , \137 , \138 , \139 , \140 , \141 , \142 , \143 , \144 , \145 ,         \146 , \147 , \148 , \149 , \150 , \151 , \152 , \153 , \154 , \155_ONE ,         \156_A[0] , \157_B[0] , \158 , \159_Z[0] , \160 , \161_A[1] , \162 , \163_B[1] , \164 , \165 ,         \166_Z[1] , \167_A[2] , \168 , \169 , \170 , \171 , \172 , \173_B[2] , \174 , \175 ,         \176_Z[2] , \177_A[3] , \178 , \179 , \180 , \181 , \182 , \183 , \184 , \185 ,         \186 , \187 , \188 , \189_B[3] , \190 , \191 , \192_Z[3] , \193_A[4] , \194 , \195 ,         \196 , \197 , \198 , \199 , \200 , \201 , \202 , \203 , \204 , \205 ,         \206 , \207 , \208 , \209 , \210 , \211_B[4] , \212 , \213 , \214_Z[4] , \215_A[5] ,         \216 , \217 , \218 , \219 , \220 , \221 , \222 , \223 , \224 , \225 ,         \226 , \227 , \228 , \229 , \230 , \231 , \232 , \233 , \234 , \235 ,         \236 , \237 , \238 , \239_B[5] , \240 , \241 , \242_Z[5] , \243_A[6] , \244 , \245 ,         \246 , \247 , \248 , \249 , \250 , \251 , \252 , \253 , \254 , \255 ,         \256 , \257 , \258 , \259 , \260 , \261 , \262 , \263 , \264 , \265 ,         \266 , \267 , \268 , \269 , \270 , \271 , \272 , \273_B[6] , \274 , \275 ,         \276_Z[6] , \277_A[7] , \278 , \279 , \280 , \281 , \282 , \283 , \284 , \285 ,         \286 , \287 , \288 , \289 , \290 , \291 , \292 , \293 , \294 , \295 ,         \296 , \297 , \298 , \299 , \300 , \301 , \302 , \303 , \304 , \305 ,         \306 , \307 , \308 , \309 , \310 , \311 , \312 , \313_B[7] , \314 , \315 ,         \316_Z[7] , \317_A[8] , \318 , \319 , \320 , \321 , \322 , \323 , \324 , \325 ,         \326 , \327 , \328 , \329 , \330 , \331 , \332 , \333 , \334 , \335 ,         \336 , \337 , \338 , \339 , \340 , \341 , \342 , \343 , \344 , \345 ,         \346 , \347 , \348 , \349 , \350 , \351 , \352 , \353 , \354 , \355 ,         \356 , \357 , \358 , \359_B[8] , \360 , \361 , \362_Z[8] , \363_A[9] , \364 , \365 ,         \366 , \367 , \368 , \369 , \370 , \371 , \372 , \373 , \374 , \375 ,         \376 , \377 , \378 , \379 , \380 , \381 , \382 , \383 , \384 , \385 ,         \386 , \387 , \388 , \389 , \390 , \391 , \392 , \393 , \394 , \395 ,         \396 , \397 , \398 , \399 , \400 , \401 , \402 , \403 , \404 , \405 ,         \406 , \407 , \408 , \409 , \410 , \411_B[9] , \412 , \413 , \414_Z[9] , \415_A[10] ,         \416 , \417 , \418 , \419 , \420 , \421 , \422 , \423 , \424 , \425 ,         \426 , \427 , \428 , \429 , \430 , \431 , \432 , \433 , \434 , \435 ,         \436 , \437 , \438 , \439 , \440 , \441 , \442 , \443 , \444 , \445 ,         \446 , \447 , \448 , \449 , \450 , \451 , \452 , \453 , \454 , \455 ,         \456 , \457 , \458 , \459 , \460 , \461 , \462 , \463 , \464 , \465 ,         \466 , \467 , \468 , \469_B[10] , \470 , \471 , \472_Z[10] , \473_A[11] , \474 , \475 ,         \476 , \477 , \478 , \479 , \480 , \481 , \482 , \483 , \484 , \485 ,         \486 , \487 , \488 , \489 , \490 , \491 , \492 , \493 , \494 , \495 ,         \496 , \497 , \498 , \499 , \500 , \501 , \502 , \503 , \504 , \505 ,         \506 , \507 , \508 , \509 , \510 , \511 , \512 , \513 , \514 , \515 ,         \516 , \517 , \518 , \519 , \520 , \521 , \522 , \523 , \524 , \525 ,         \526 , \527 , \528 , \529 , \530 , \531 , \532 , \533_B[11] , \534 , \535 ,         \536_Z[11] , \537_A[12] , \538 , \539 , \540 , \541 , \542 , \543 , \544 , \545 ,         \546 , \547 , \548 , \549 , \550 , \551 , \552 , \553 , \554 , \555 ,         \556 , \557 , \558 , \559 , \560 , \561 , \562 , \563 , \564 , \565 ,         \566 , \567 , \568 , \569 , \570 , \571 , \572 , \573 , \574 , \575 ,         \576 , \577 , \578 , \579 , \580 , \581 , \582 , \583 , \584 , \585 ,         \586 , \587 , \588 , \589 , \590 , \591 , \592 , \593 , \594 , \595 ,         \596 , \597 , \598 , \599 , \600 , \601 , \602 , \603_B[12] , \604 , \605 ,         \606_Z[12] , \607_A[13] , \608 , \609 , \610 , \611 , \612 , \613 , \614 , \615 ,         \616 , \617 , \618 , \619 , \620 , \621 , \622 , \623 , \624 , \625 ,         \626 , \627 , \628 , \629 , \630 , \631 , \632 , \633 , \634 , \635 ,         \636 , \637 , \638 , \639 , \640 , \641 , \642 , \643 , \644 , \645 ,         \646 , \647 , \648 , \649 , \650 , \651 , \652 , \653 , \654 , \655 ,         \656 , \657 , \658 , \659 , \660 , \661 , \662 , \663 , \664 , \665 ,         \666 , \667 , \668 , \669 , \670 , \671 , \672 , \673 , \674 , \675 ,         \676 , \677 , \678 , \679_B[13] , \680 , \681 , \682_Z[13] , \683_A[14] , \684 , \685 ,         \686 , \687 , \688 , \689 , \690 , \691 , \692 , \693 , \694 , \695 ,         \696 , \697 , \698 , \699 , \700 , \701 , \702 , \703 , \704 , \705 ,         \706 , \707 , \708 , \709 , \710 , \711 , \712 , \713 , \714 , \715 ,         \716 , \717 , \718 , \719 , \720 , \721 , \722 , \723 , \724 , \725 ,         \726 , \727 , \728 , \729 , \730 , \731 , \732 , \733 , \734 , \735 ,         \736 , \737 , \738 , \739 , \740 , \741 , \742 , \743 , \744 , \745 ,         \746 , \747 , \748 , \749 , \750 , \751 , \752 , \753 , \754 , \755 ,         \756 , \757 , \758 , \759 , \760 , \761_B[14] , \762 , \763 , \764_Z[14] , \765_A[15] ,         \766 , \767 , \768 , \769 , \770 , \771 , \772 , \773 , \774 , \775 ,         \776 , \777 , \778 , \779 , \780 , \781 , \782 , \783 , \784 , \785 ,         \786 , \787 , \788 , \789 , \790 , \791 , \792 , \793 , \794 , \795 ,         \796 , \797 , \798 , \799 , \800 , \801 , \802 , \803 , \804 , \805 ,         \806 , \807 , \808 , \809 , \810 , \811 , \812 , \813 , \814 , \815 ,         \816 , \817 , \818 , \819 , \820 , \821 , \822 , \823 , \824 , \825 ,         \826 , \827 , \828 , \829 , \830 , \831 , \832 , \833 , \834 , \835 ,         \836 , \837 , \838 , \839 , \840 , \841 , \842 , \843 , \844 , \845 ,         \846 , \847 , \848 , \849_B[15] , \850 , \851 , \852_Z[15] , \853 , \854 , \855 ,         \856 , \857 , \858 , \859 , \860 , \861 , \862 , \863 , \864 , \865 ,         \866 , \867 , \868 , \869 , \870 , \871 , \872 , \873 , \874 , \875 ,         \876 , \877 , \878 , \879 , \880 , \881 , \882 , \883 , \884 , \885 ,         \886_A[0] , \887_B[0] , \888 , \889_Z[0] , \890 , \891_A[0] , \892_B[0] , \893 , \894_Z[0] , \895 ,         \896_A[0] , \897_B[0] , \898 , \899_SUM[0] , \900 , \901_A[0] , \902_B[0] , \903 , \904_SUM[0] , \905 ,         \906 , \907 , \908 , \909 , \910 , \911 , \912 , \913 , \914 , \915 ,         \916 , \917 , \918 , \919 , \920_A[1] , \921 , \922_B[1] , \923 , \924 , \925_Z[1] ,         \926 , \927_A[1] , \928 , \929_B[1] , \930 , \931 , \932_Z[1] , \933 , \934_A[1] , \935_B[1] ,         \936 , \937 , \938 , \939_SUM[1] , \940 , \941_A[1] , \942_B[1] , \943 , \944 , \945 ,         \946_SUM[1] , \947 , \948 , \949 , \950 , \951 , \952 , \953 , \954 , \955 ,         \956 , \957 , \958 , \959 , \960 , \961 , \962_A[2] , \963 , \964 , \965 ,         \966 , \967 , \968_B[2] , \969 , \970 , \971_Z[2] , \972 , \973_A[2] , \974 , \975 ,         \976 , \977 , \978 , \979_B[2] , \980 , \981 , \982_Z[2] , \983 , \984_A[2] , \985_B[2] ,         \986 , \987 , \988 , \989 , \990 , \991 , \992_SUM[2] , \993 , \994_A[2] , \995_B[2] ,         \996 , \997 , \998 , \999 , \1000 , \1001 , \1002_SUM[2] , \1003 , \1004 , \1005 ,         \1006 , \1007 , \1008 , \1009 , \1010 , \1011 , \1012 , \1013 , \1014 , \1015 ,         \1016 , \1017 , \1018_A[3] , \1019 , \1020 , \1021 , \1022 , \1023 , \1024 , \1025 ,         \1026 , \1027 , \1028 , \1029 , \1030_B[3] , \1031 , \1032 , \1033_Z[3] , \1034 , \1035_A[3] ,         \1036 , \1037 , \1038 , \1039 , \1040 , \1041 , \1042 , \1043 , \1044 , \1045 ,         \1046 , \1047_B[3] , \1048 , \1049 , \1050_Z[3] , \1051 , \1052_A[3] , \1053_B[3] , \1054 , \1055 ,         \1056 , \1057 , \1058 , \1059 , \1060_SUM[3] , \1061 , \1062_A[3] , \1063_B[3] , \1064 , \1065 ,         \1066 , \1067 , \1068 , \1069 , \1070_SUM[3] , \1071 , \1072 , \1073 , \1074 , \1075 ,         \1076 , \1077 , \1078 , \1079 , \1080 , \1081 , \1082 , \1083 , \1084 , \1085 ,         \1086_A[4] , \1087 , \1088 , \1089 , \1090 , \1091 , \1092 , \1093 , \1094 , \1095 ,         \1096 , \1097 , \1098 , \1099 , \1100 , \1101 , \1102 , \1103 , \1104_B[4] , \1105 ,         \1106 , \1107_Z[4] , \1108 , \1109_A[4] , \1110 , \1111 , \1112 , \1113 , \1114 , \1115 ,         \1116 , \1117 , \1118 , \1119 , \1120 , \1121 , \1122 , \1123 , \1124 , \1125 ,         \1126 , \1127_B[4] , \1128 , \1129 , \1130_Z[4] , \1131 , \1132_A[4] , \1133_B[4] , \1134 , \1135 ,         \1136 , \1137 , \1138 , \1139 , \1140_SUM[4] , \1141 , \1142_A[4] , \1143_B[4] , \1144 , \1145 ,         \1146 , \1147 , \1148 , \1149 , \1150_SUM[4] , \1151 , \1152 , \1153 , \1154 , \1155 ,         \1156 , \1157 , \1158 , \1159 , \1160 , \1161 , \1162 , \1163 , \1164 , \1165 ,         \1166_A[5] , \1167 , \1168 , \1169 , \1170 , \1171 , \1172 , \1173 , \1174 , \1175 ,         \1176 , \1177 , \1178 , \1179 , \1180 , \1181 , \1182 , \1183 , \1184 , \1185 ,         \1186 , \1187 , \1188 , \1189 , \1190_B[5] , \1191 , \1192 , \1193_Z[5] , \1194 , \1195_A[5] ,         \1196 , \1197 , \1198 , \1199 , \1200 , \1201 , \1202 , \1203 , \1204 , \1205 ,         \1206 , \1207 , \1208 , \1209 , \1210 , \1211 , \1212 , \1213 , \1214 , \1215 ,         \1216 , \1217 , \1218 , \1219_B[5] , \1220 , \1221 , \1222_Z[5] , \1223 , \1224_A[5] , \1225_B[5] ,         \1226 , \1227 , \1228 , \1229 , \1230 , \1231 , \1232_SUM[5] , \1233 , \1234_A[5] , \1235_B[5] ,         \1236 , \1237 , \1238 , \1239 , \1240 , \1241 , \1242_SUM[5] , \1243 , \1244 , \1245 ,         \1246 , \1247 , \1248 , \1249 , \1250 , \1251 , \1252 , \1253 , \1254 , \1255 ,         \1256 , \1257 , \1258_A[6] , \1259 , \1260 , \1261 , \1262 , \1263 , \1264 , \1265 ,         \1266 , \1267 , \1268 , \1269 , \1270 , \1271 , \1272 , \1273 , \1274 , \1275 ,         \1276 , \1277 , \1278 , \1279 , \1280 , \1281 , \1282 , \1283 , \1284 , \1285 ,         \1286 , \1287 , \1288_B[6] , \1289 , \1290 , \1291_Z[6] , \1292 , \1293_A[6] , \1294 , \1295 ,         \1296 , \1297 , \1298 , \1299 , \1300 , \1301 , \1302 , \1303 , \1304 , \1305 ,         \1306 , \1307 , \1308 , \1309 , \1310 , \1311 , \1312 , \1313 , \1314 , \1315 ,         \1316 , \1317 , \1318 , \1319 , \1320 , \1321 , \1322 , \1323_B[6] , \1324 , \1325 ,         \1326_Z[6] , \1327 , \1328_A[6] , \1329_B[6] , \1330 , \1331 , \1332 , \1333 , \1334 , \1335 ,         \1336_SUM[6] , \1337 , \1338_A[6] , \1339_B[6] , \1340 , \1341 , \1342 , \1343 , \1344 , \1345 ,         \1346_SUM[6] , \1347 , \1348 , \1349 , \1350 , \1351 , \1352 , \1353 , \1354 , \1355 ,         \1356 , \1357 , \1358 , \1359 , \1360 , \1361 , \1362_A[7] , \1363 , \1364 , \1365 ,         \1366 , \1367 , \1368 , \1369 , \1370 , \1371 , \1372 , \1373 , \1374 , \1375 ,         \1376 , \1377 , \1378 , \1379 , \1380 , \1381 , \1382 , \1383 , \1384 , \1385 ,         \1386 , \1387 , \1388 , \1389 , \1390 , \1391 , \1392 , \1393 , \1394 , \1395 ,         \1396 , \1397 , \1398_B[7] , \1399 , \1400 , \1401_Z[7] , \1402 , \1403_A[7] , \1404 , \1405 ,         \1406 , \1407 , \1408 , \1409 , \1410 , \1411 , \1412 , \1413 , \1414 , \1415 ,         \1416 , \1417 , \1418 , \1419 , \1420 , \1421 , \1422 , \1423 , \1424 , \1425 ,         \1426 , \1427 , \1428 , \1429 , \1430 , \1431 , \1432 , \1433 , \1434 , \1435 ,         \1436 , \1437 , \1438 , \1439_B[7] , \1440 , \1441 , \1442_Z[7] , \1443 , \1444_A[7] , \1445_B[7] ,         \1446 , \1447 , \1448 , \1449 , \1450 , \1451 , \1452_SUM[7] , \1453 , \1454_A[7] , \1455_B[7] ,         \1456 , \1457 , \1458 , \1459 , \1460 , \1461 , \1462_SUM[7] , \1463 , \1464 , \1465 ,         \1466 , \1467 , \1468 , \1469 , \1470 , \1471 , \1472 , \1473 , \1474 , \1475 ,         \1476 , \1477 , \1478_A[8] , \1479 , \1480 , \1481 , \1482 , \1483 , \1484 , \1485 ,         \1486 , \1487 , \1488 , \1489 , \1490 , \1491 , \1492 , \1493 , \1494 , \1495 ,         \1496 , \1497 , \1498 , \1499 , \1500 , \1501 , \1502 , \1503 , \1504 , \1505 ,         \1506 , \1507 , \1508 , \1509 , \1510 , \1511 , \1512 , \1513 , \1514 , \1515 ,         \1516 , \1517 , \1518 , \1519 , \1520_B[8] , \1521 , \1522 , \1523_Z[8] , \1524 , \1525_A[8] ,         \1526 , \1527 , \1528 , \1529 , \1530 , \1531 , \1532 , \1533 , \1534 , \1535 ,         \1536 , \1537 , \1538 , \1539 , \1540 , \1541 , \1542 , \1543 , \1544 , \1545 ,         \1546 , \1547 , \1548 , \1549 , \1550 , \1551 , \1552 , \1553 , \1554 , \1555 ,         \1556 , \1557 , \1558 , \1559 , \1560 , \1561 , \1562 , \1563 , \1564 , \1565 ,         \1566 , \1567_B[8] , \1568 , \1569 , \1570_Z[8] , \1571 , \1572_A[8] , \1573_B[8] , \1574 , \1575 ,         \1576 , \1577 , \1578 , \1579 , \1580_SUM[8] , \1581 , \1582_A[8] , \1583_B[8] , \1584 , \1585 ,         \1586 , \1587 , \1588 , \1589 , \1590_SUM[8] , \1591 , \1592 , \1593 , \1594 , \1595 ,         \1596 , \1597 , \1598 , \1599 , \1600 , \1601 , \1602 , \1603 , \1604 , \1605 ,         \1606_A[9] , \1607 , \1608 , \1609 , \1610 , \1611 , \1612 , \1613 , \1614 , \1615 ,         \1616 , \1617 , \1618 , \1619 , \1620 , \1621 , \1622 , \1623 , \1624 , \1625 ,         \1626 , \1627 , \1628 , \1629 , \1630 , \1631 , \1632 , \1633 , \1634 , \1635 ,         \1636 , \1637 , \1638 , \1639 , \1640 , \1641 , \1642 , \1643 , \1644 , \1645 ,         \1646 , \1647 , \1648 , \1649 , \1650 , \1651 , \1652 , \1653 , \1654_B[9] , \1655 ,         \1656 , \1657_Z[9] , \1658 , \1659_A[9] , \1660 , \1661 , \1662 , \1663 , \1664 , \1665 ,         \1666 , \1667 , \1668 , \1669 , \1670 , \1671 , \1672 , \1673 , \1674 , \1675 ,         \1676 , \1677 , \1678 , \1679 , \1680 , \1681 , \1682 , \1683 , \1684 , \1685 ,         \1686 , \1687 , \1688 , \1689 , \1690 , \1691 , \1692 , \1693 , \1694 , \1695 ,         \1696 , \1697 , \1698 , \1699 , \1700 , \1701 , \1702 , \1703 , \1704 , \1705 ,         \1706 , \1707_B[9] , \1708 , \1709 , \1710_Z[9] , \1711 , \1712_A[9] , \1713_B[9] , \1714 , \1715 ,         \1716 , \1717 , \1718 , \1719 , \1720_SUM[9] , \1721 , \1722_A[9] , \1723_B[9] , \1724 , \1725 ,         \1726 , \1727 , \1728 , \1729 , \1730_SUM[9] , \1731 , \1732 , \1733 , \1734 , \1735 ,         \1736 , \1737 , \1738 , \1739 , \1740 , \1741 , \1742 , \1743 , \1744 , \1745 ,         \1746_A[10] , \1747 , \1748 , \1749 , \1750 , \1751 , \1752 , \1753 , \1754 , \1755 ,         \1756 , \1757 , \1758 , \1759 , \1760 , \1761 , \1762 , \1763 , \1764 , \1765 ,         \1766 , \1767 , \1768 , \1769 , \1770 , \1771 , \1772 , \1773 , \1774 , \1775 ,         \1776 , \1777 , \1778 , \1779 , \1780 , \1781 , \1782 , \1783 , \1784 , \1785 ,         \1786 , \1787 , \1788 , \1789 , \1790 , \1791 , \1792 , \1793 , \1794 , \1795 ,         \1796 , \1797 , \1798 , \1799 , \1800_B[10] , \1801 , \1802 , \1803_Z[10] , \1804 , \1805_A[10] ,         \1806 , \1807 , \1808 , \1809 , \1810 , \1811 , \1812 , \1813 , \1814 , \1815 ,         \1816 , \1817 , \1818 , \1819 , \1820 , \1821 , \1822 , \1823 , \1824 , \1825 ,         \1826 , \1827 , \1828 , \1829 , \1830 , \1831 , \1832 , \1833 , \1834 , \1835 ,         \1836 , \1837 , \1838 , \1839 , \1840 , \1841 , \1842 , \1843 , \1844 , \1845 ,         \1846 , \1847 , \1848 , \1849 , \1850 , \1851 , \1852 , \1853 , \1854 , \1855 ,         \1856 , \1857 , \1858 , \1859_B[10] , \1860 , \1861 , \1862_Z[10] , \1863 , \1864_A[10] , \1865_B[10] ,         \1866 , \1867 , \1868 , \1869 , \1870 , \1871 , \1872_SUM[10] , \1873 , \1874_A[10] , \1875_B[10] ,         \1876 , \1877 , \1878 , \1879 , \1880 , \1881 , \1882_SUM[10] , \1883 , \1884 , \1885 ,         \1886 , \1887 , \1888 , \1889 , \1890 , \1891 , \1892 , \1893 , \1894 , \1895 ,         \1896 , \1897 , \1898_A[11] , \1899 , \1900 , \1901 , \1902 , \1903 , \1904 , \1905 ,         \1906 , \1907 , \1908 , \1909 , \1910 , \1911 , \1912 , \1913 , \1914 , \1915 ,         \1916 , \1917 , \1918 , \1919 , \1920 , \1921 , \1922 , \1923 , \1924 , \1925 ,         \1926 , \1927 , \1928 , \1929 , \1930 , \1931 , \1932 , \1933 , \1934 , \1935 ,         \1936 , \1937 , \1938 , \1939 , \1940 , \1941 , \1942 , \1943 , \1944 , \1945 ,         \1946 , \1947 , \1948 , \1949 , \1950 , \1951 , \1952 , \1953 , \1954 , \1955 ,         \1956 , \1957 , \1958_B[11] , \1959 , \1960 , \1961_Z[11] , \1962 , \1963_A[11] , \1964 , \1965 ,         \1966 , \1967 , \1968 , \1969 , \1970 , \1971 , \1972 , \1973 , \1974 , \1975 ,         \1976 , \1977 , \1978 , \1979 , \1980 , \1981 , \1982 , \1983 , \1984 , \1985 ,         \1986 , \1987 , \1988 , \1989 , \1990 , \1991 , \1992 , \1993 , \1994 , \1995 ,         \1996 , \1997 , \1998 , \1999 , \2000 , \2001 , \2002 , \2003 , \2004 , \2005 ,         \2006 , \2007 , \2008 , \2009 , \2010 , \2011 , \2012 , \2013 , \2014 , \2015 ,         \2016 , \2017 , \2018 , \2019 , \2020 , \2021 , \2022 , \2023_B[11] , \2024 , \2025 ,         \2026_Z[11] , \2027 , \2028_A[11] , \2029_B[11] , \2030 , \2031 , \2032 , \2033 , \2034 , \2035 ,         \2036_SUM[11] , \2037 , \2038_A[11] , \2039_B[11] , \2040 , \2041 , \2042 , \2043 , \2044 , \2045 ,         \2046_SUM[11] , \2047 , \2048 , \2049 , \2050 , \2051 , \2052 , \2053 , \2054 , \2055 ,         \2056 , \2057 , \2058 , \2059 , \2060 , \2061 , \2062_A[12] , \2063 , \2064 , \2065 ,         \2066 , \2067 , \2068 , \2069 , \2070 , \2071 , \2072 , \2073 , \2074 , \2075 ,         \2076 , \2077 , \2078 , \2079 , \2080 , \2081 , \2082 , \2083 , \2084 , \2085 ,         \2086 , \2087 , \2088 , \2089 , \2090 , \2091 , \2092 , \2093 , \2094 , \2095 ,         \2096 , \2097 , \2098 , \2099 , \2100 , \2101 , \2102 , \2103 , \2104 , \2105 ,         \2106 , \2107 , \2108 , \2109 , \2110 , \2111 , \2112 , \2113 , \2114 , \2115 ,         \2116 , \2117 , \2118 , \2119 , \2120 , \2121 , \2122 , \2123 , \2124 , \2125 ,         \2126 , \2127 , \2128_B[12] , \2129 , \2130 , \2131_Z[12] , \2132 , \2133_A[12] , \2134 , \2135 ,         \2136 , \2137 , \2138 , \2139 , \2140 , \2141 , \2142 , \2143 , \2144 , \2145 ,         \2146 , \2147 , \2148 , \2149 , \2150 , \2151 , \2152 , \2153 , \2154 , \2155 ,         \2156 , \2157 , \2158 , \2159 , \2160 , \2161 , \2162 , \2163 , \2164 , \2165 ,         \2166 , \2167 , \2168 , \2169 , \2170 , \2171 , \2172 , \2173 , \2174 , \2175 ,         \2176 , \2177 , \2178 , \2179 , \2180 , \2181 , \2182 , \2183 , \2184 , \2185 ,         \2186 , \2187 , \2188 , \2189 , \2190 , \2191 , \2192 , \2193 , \2194 , \2195 ,         \2196 , \2197 , \2198 , \2199_B[12] , \2200 , \2201 , \2202_Z[12] , \2203 , \2204_A[12] , \2205_B[12] ,         \2206 , \2207 , \2208 , \2209 , \2210 , \2211 , \2212_SUM[12] , \2213 , \2214_A[12] , \2215_B[12] ,         \2216 , \2217 , \2218 , \2219 , \2220 , \2221 , \2222_SUM[12] , \2223 , \2224 , \2225 ,         \2226 , \2227 , \2228 , \2229 , \2230 , \2231 , \2232 , \2233 , \2234 , \2235 ,         \2236 , \2237 , \2238_A[13] , \2239 , \2240 , \2241 , \2242 , \2243 , \2244 , \2245 ,         \2246 , \2247 , \2248 , \2249 , \2250 , \2251 , \2252 , \2253 , \2254 , \2255 ,         \2256 , \2257 , \2258 , \2259 , \2260 , \2261 , \2262 , \2263 , \2264 , \2265 ,         \2266 , \2267 , \2268 , \2269 , \2270 , \2271 , \2272 , \2273 , \2274 , \2275 ,         \2276 , \2277 , \2278 , \2279 , \2280 , \2281 , \2282 , \2283 , \2284 , \2285 ,         \2286 , \2287 , \2288 , \2289 , \2290 , \2291 , \2292 , \2293 , \2294 , \2295 ,         \2296 , \2297 , \2298 , \2299 , \2300 , \2301 , \2302 , \2303 , \2304 , \2305 ,         \2306 , \2307 , \2308 , \2309 , \2310_B[13] , \2311 , \2312 , \2313_Z[13] , \2314 , \2315_A[13] ,         \2316 , \2317 , \2318 , \2319 , \2320 , \2321 , \2322 , \2323 , \2324 , \2325 ,         \2326 , \2327 , \2328 , \2329 , \2330 , \2331 , \2332 , \2333 , \2334 , \2335 ,         \2336 , \2337 , \2338 , \2339 , \2340 , \2341 , \2342 , \2343 , \2344 , \2345 ,         \2346 , \2347 , \2348 , \2349 , \2350 , \2351 , \2352 , \2353 , \2354 , \2355 ,         \2356 , \2357 , \2358 , \2359 , \2360 , \2361 , \2362 , \2363 , \2364 , \2365 ,         \2366 , \2367 , \2368 , \2369 , \2370 , \2371 , \2372 , \2373 , \2374 , \2375 ,         \2376 , \2377 , \2378 , \2379 , \2380 , \2381 , \2382 , \2383 , \2384 , \2385 ,         \2386 , \2387_B[13] , \2388 , \2389 , \2390_Z[13] , \2391 , \2392_A[13] , \2393_B[13] , \2394 , \2395 ,         \2396 , \2397 , \2398 , \2399 , \2400_SUM[13] , \2401 , \2402_A[13] , \2403_B[13] , \2404 , \2405 ,         \2406 , \2407 , \2408 , \2409 , \2410_SUM[13] , \2411 , \2412 , \2413 , \2414 , \2415 ,         \2416 , \2417 , \2418 , \2419 , \2420 , \2421 , \2422 , \2423 , \2424 , \2425 ,         \2426_A[14] , \2427 , \2428 , \2429 , \2430 , \2431 , \2432 , \2433 , \2434 , \2435 ,         \2436 , \2437 , \2438 , \2439 , \2440 , \2441 , \2442 , \2443 , \2444 , \2445 ,         \2446 , \2447 , \2448 , \2449 , \2450 , \2451 , \2452 , \2453 , \2454 , \2455 ,         \2456 , \2457 , \2458 , \2459 , \2460 , \2461 , \2462 , \2463 , \2464 , \2465 ,         \2466 , \2467 , \2468 , \2469 , \2470 , \2471 , \2472 , \2473 , \2474 , \2475 ,         \2476 , \2477 , \2478 , \2479 , \2480 , \2481 , \2482 , \2483 , \2484 , \2485 ,         \2486 , \2487 , \2488 , \2489 , \2490 , \2491 , \2492 , \2493 , \2494 , \2495 ,         \2496 , \2497 , \2498 , \2499 , \2500 , \2501 , \2502 , \2503 , \2504_B[14] , \2505 ,         \2506 , \2507_Z[14] , \2508 , \2509_A[14] , \2510 , \2511 , \2512 , \2513 , \2514 , \2515 ,         \2516 , \2517 , \2518 , \2519 , \2520 , \2521 , \2522 , \2523 , \2524 , \2525 ,         \2526 , \2527 , \2528 , \2529 , \2530 , \2531 , \2532 , \2533 , \2534 , \2535 ,         \2536 , \2537 , \2538 , \2539 , \2540 , \2541 , \2542 , \2543 , \2544 , \2545 ,         \2546 , \2547 , \2548 , \2549 , \2550 , \2551 , \2552 , \2553 , \2554 , \2555 ,         \2556 , \2557 , \2558 , \2559 , \2560 , \2561 , \2562 , \2563 , \2564 , \2565 ,         \2566 , \2567 , \2568 , \2569 , \2570 , \2571 , \2572 , \2573 , \2574 , \2575 ,         \2576 , \2577 , \2578 , \2579 , \2580 , \2581 , \2582 , \2583 , \2584 , \2585 ,         \2586 , \2587_B[14] , \2588 , \2589 , \2590_Z[14] , \2591 , \2592_A[14] , \2593_B[14] , \2594 , \2595 ,         \2596 , \2597 , \2598 , \2599 , \2600_SUM[14] , \2601 , \2602_A[14] , \2603_B[14] , \2604 , \2605 ,         \2606 , \2607 , \2608 , \2609 , \2610_SUM[14] , \2611 , \2612 , \2613 , \2614 , \2615 ,         \2616 , \2617 , \2618 , \2619 , \2620 , \2621 , \2622 , \2623 , \2624 , \2625 ,         \2626_A[15] , \2627 , \2628 , \2629 , \2630 , \2631 , \2632 , \2633 , \2634 , \2635 ,         \2636 , \2637 , \2638 , \2639 , \2640 , \2641 , \2642 , \2643 , \2644 , \2645 ,         \2646 , \2647 , \2648 , \2649 , \2650 , \2651 , \2652 , \2653 , \2654 , \2655 ,         \2656 , \2657 , \2658 , \2659 , \2660 , \2661 , \2662 , \2663 , \2664 , \2665 ,         \2666 , \2667 , \2668 , \2669 , \2670 , \2671 , \2672 , \2673 , \2674 , \2675 ,         \2676 , \2677 , \2678 , \2679 , \2680 , \2681 , \2682 , \2683 , \2684 , \2685 ,         \2686 , \2687 , \2688 , \2689 , \2690 , \2691 , \2692 , \2693 , \2694 , \2695 ,         \2696 , \2697 , \2698 , \2699 , \2700 , \2701 , \2702 , \2703 , \2704 , \2705 ,         \2706 , \2707 , \2708 , \2709 , \2710_B[15] , \2711 , \2712 , \2713_Z[15] , \2714 , \2715_A[15] ,         \2716 , \2717 , \2718 , \2719 , \2720 , \2721 , \2722 , \2723 , \2724 , \2725 ,         \2726 , \2727 , \2728 , \2729 , \2730 , \2731 , \2732 , \2733 , \2734 , \2735 ,         \2736 , \2737 , \2738 , \2739 , \2740 , \2741 , \2742 , \2743 , \2744 , \2745 ,         \2746 , \2747 , \2748 , \2749 , \2750 , \2751 , \2752 , \2753 , \2754 , \2755 ,         \2756 , \2757 , \2758 , \2759 , \2760 , \2761 , \2762 , \2763 , \2764 , \2765 ,         \2766 , \2767 , \2768 , \2769 , \2770 , \2771 , \2772 , \2773 , \2774 , \2775 ,         \2776 , \2777 , \2778 , \2779 , \2780 , \2781 , \2782 , \2783 , \2784 , \2785 ,         \2786 , \2787 , \2788 , \2789 , \2790 , \2791 , \2792 , \2793 , \2794 , \2795 ,         \2796 , \2797 , \2798 , \2799_B[15] , \2800 , \2801 , \2802_Z[15] , \2803 , \2804_A[15] , \2805_B[15] ,         \2806 , \2807 , \2808 , \2809 , \2810 , \2811 , \2812_SUM[15] , \2813 , \2814_A[15] , \2815_B[15] ,         \2816 , \2817 , \2818 , \2819 , \2820 , \2821 , \2822_SUM[15] , \2823 , \2824 , \2825 ,         \2826 , \2827 , \2828 , \2829_A[15] , \2830_B[15] , \2831 , \2832_A[14] , \2833_B[14] , \2834 , \2835_A[13] ,         \2836_B[13] , \2837 , \2838_A[12] , \2839_B[12] , \2840 , \2841_A[11] , \2842_B[11] , \2843 , \2844_A[10] , \2845_B[10] ,         \2846 , \2847_A[9] , \2848_B[9] , \2849 , \2850_A[8] , \2851_B[8] , \2852 , \2853_A[7] , \2854_B[7] , \2855 ,         \2856_A[6] , \2857_B[6] , \2858 , \2859_A[5] , \2860_B[5] , \2861 , \2862_A[4] , \2863_B[4] , \2864 , \2865_A[3] ,         \2866_B[3] , \2867 , \2868_A[2] , \2869_B[2] , \2870 , \2871_A[1] , \2872_B[1] , \2873 , \2874_A[0] , \2875_B[0] ,         \2876 , \2877 , \2878 , \2879 , \2880 , \2881 , \2882 , \2883 , \2884 , \2885 ,         \2886 , \2887 , \2888 , \2889 , \2890 , \2891 , \2892 , \2893 , \2894 , \2895 ,         \2896 , \2897 , \2898 , \2899 , \2900 , \2901 , \2902 , \2903 , \2904 , \2905 ,         \2906 , \2907 , \2908 , \2909 , \2910 , \2911 , \2912 , \2913 , \2914 , \2915 ,         \2916 , \2917 , \2918 , \2919 , \2920 , \2921 , \2922_SUM[16] , \2923_A[16] , \2924 , \2925 ,         \2926_SUM[15] , \2927_A[15] , \2928 , \2929 , \2930_SUM[14] , \2931_A[14] , \2932 , \2933 , \2934_SUM[13] , \2935_A[13] ,         \2936 , \2937 , \2938_SUM[12] , \2939_A[12] , \2940 , \2941 , \2942_SUM[11] , \2943_A[11] , \2944 , \2945 ,         \2946_SUM[10] , \2947_A[10] , \2948 , \2949 , \2950_SUM[9] , \2951_A[9] , \2952 , \2953 , \2954_SUM[8] , \2955_A[8] ,         \2956 , \2957 , \2958_SUM[7] , \2959_A[7] , \2960 , \2961 , \2962_SUM[6] , \2963_A[6] , \2964 , \2965 ,         \2966_SUM[5] , \2967_A[5] , \2968 , \2969 , \2970_SUM[4] , \2971_A[4] , \2972 , \2973 , \2974_SUM[3] , \2975_A[3] ,         \2976 , \2977 , \2978_SUM[2] , \2979_A[2] , \2980 , \2981 , \2982_SUM[1] , \2983_A[1] , \2984 , \2985_SUM[0] ,         \2986_A[0] , \2987_B[15] , \2988_B[14] , \2989_B[13] , \2990_B[12] , \2991_B[11] , \2992_B[10] , \2993_B[9] , \2994_B[8] , \2995_B[7] ,         \2996_B[6] , \2997_B[5] , \2998_B[4] , \2999_B[3] , \3000_B[2] , \3001_B[1] , \3002_B[0] , \3003 , \3004 , \3005 ,         \3006 , \3007 , \3008 , \3009 , \3010 , \3011 , \3012 , \3013 , \3014 , \3015 ,         \3016 , \3017 , \3018 , \3019 , \3020 , \3021 , \3022 , \3023 , \3024 , \3025 ,         \3026 , \3027 , \3028 , \3029 , \3030 , \3031 , \3032 , \3033 , \3034 , \3035 ,         \3036 , \3037 , \3038 , \3039 , \3040 , \3041 , \3042 , \3043 , \3044 , \3045 ,         \3046 , \3047 , \3048 , \3049 , \3050 , \3051 , \3052 , \3053 , \3054 , \3055 ,         \3056 , \3057 , \3058 , \3059 , \3060 , \3061 , \3062 , \3063 , \3064 , \3065 ,         \3066 , \3067 , \3068 , \3069 , \3070 , \3071 , \3072 , \3073 , \3074 , \3075 ,         \3076 , \3077 , \3078 , \3079 , \3080 , \3081 , \3082 , \3083 , \3084 , \3085 ,         \3086 , \3087 , \3088 , \3089 , \3090 , \3091 , \3092 , \3093 , \3094 , \3095 ,         \3096 , \3097 , \3098 , \3099 , \3100 , \3101 , \3102 , \3103 , \3104 , \3105 ,         \3106 , \3107 , \3108 , \3109 , \3110 , \3111 , \3112 , \3113 , \3114 , \3115 ,         \3116 , \3117 , \3118 , \3119 , \3120 , \3121 , \3122 , \3123 , \3124 , \3125 ,         \3126 , \3127 , \3128 , \3129 , \3130 , \3131 , \3132 , \3133 , \3134 , \3135 ,         \3136 , \3137 , \3138 , \3139 , \3140 , \3141 , \3142 , \3143 , \3144 , \3145 ,         \3146 , \3147 , \3148 , \3149 , \3150 , \3151 , \3152 , \3153 , \3154 , \3155 ,         \3156 , \3157 , \3158 , \3159 , \3160 , \3161 , \3162 , \3163 , \3164 , \3165 ,         \3166 , \3167 , \3168 , \3169 , \3170 , \3171 , \3172 , \3173 , \3174 , \3175 ,         \3176 , \3177 , \3178 , \3179 , \3180 , \3181 , \3182 , \3183 , \3184 , \3185 ,         \3186 , \3187 , \3188 , \3189 , \3190 , \3191 , \3192 , \3193 , \3194 , \3195 ,         \3196 , \3197 , \3198 , \3199 , \3200 , \3201 , \3202 , \3203 , \3204 , \3205 ,         \3206 , \3207 , \3208 , \3209 , \3210 , \3211 , \3212 , \3213 , \3214 , \3215 ,         \3216 , \3217 , \3218 , \3219 , \3220 , \3221 , \3222 , \3223 , \3224 , \3225 ,         \3226 , \3227 , \3228 , \3229 , \3230 , \3231 , \3232 , \3233 , \3234 , \3235 ,         \3236 , \3237 , \3238 , \3239 , \3240 , \3241 , \3242 , \3243 , \3244 , \3245 ,         \3246 , \3247 , \3248 , \3249 , \3250 , \3251 , \3252 , \3253 , \3254 , \3255 ,         \3256 , \3257 , \3258 , \3259 , \3260 , \3261 , \3262 , \3263 , \3264 , \3265 ,         \3266 , \3267 , \3268 , \3269 , \3270 , \3271 , \3272 , \3273 , \3274 , \3275 ,         \3276 , \3277 , \3278 , \3279 , \3280 , \3281 , \3282 , \3283 , \3284 , \3285 ,         \3286 , \3287 , \3288 , \3289 , \3290 , \3291 , \3292 , \3293 , \3294 , \3295 ,         \3296 , \3297 , \3298 , \3299 , \3300 , \3301 , \3302 , \3303 , \3304 , \3305 ,         \3306 , \3307 , \3308 , \3309 , \3310 , \3311 , \3312 , \3313 , \3314 , \3315 ,         \3316 , \3317 , \3318 , \3319 , \3320 , \3321 , \3322 , \3323 , \3324 , \3325 ,         \3326 , \3327 , \3328 , \3329 , \3330 , \3331 , \3332 , \3333 , \3334 , \3335 ,         \3336 , \3337 , \3338 , \3339 , \3340 , \3341 , \3342 , \3343 , \3344 , \3345 ,         \3346 , \3347 , \3348 , \3349 , \3350 , \3351 , \3352 , \3353 , \3354 , \3355 ,         \3356 , \3357 , \3358 , \3359 , \3360 , \3361 , \3362 , \3363 , \3364 , \3365 ,         \3366 , \3367 , \3368 , \3369 , \3370 , \3371 , \3372 , \3373 , \3374 , \3375 ,         \3376 , \3377 , \3378 , \3379 , \3380 , \3381 , \3382 , \3383 , \3384 , \3385 ,         \3386 , \3387 , \3388 , \3389 , \3390 , \3391 , \3392 , \3393 , \3394 , \3395 ,         \3396 , \3397 , \3398 , \3399 , \3400 , \3401 , \3402 , \3403 , \3404 , \3405 ,         \3406 , \3407 , \3408 , \3409 , \3410 , \3411 , \3412 , \3413 , \3414 , \3415 ,         \3416 , \3417 , \3418 , \3419 , \3420 , \3421 , \3422 , \3423 , \3424 , \3425 ,         \3426 , \3427 , \3428 , \3429 , \3430 , \3431 , \3432 , \3433 , \3434 , \3435 ,         \3436 , \3437 , \3438 , \3439 , \3440 , \3441 , \3442 , \3443 , \3444 , \3445 ,         \3446 , \3447 , \3448 , \3449 , \3450 , \3451 , \3452 , \3453 , \3454 , \3455 ,         \3456 , \3457 , \3458 , \3459 , \3460 , \3461 , \3462 , \3463 , \3464 , \3465 ,         \3466 , \3467 , \3468 , \3469 , \3470 , \3471 , \3472 , \3473 , \3474 , \3475 ,         \3476 , \3477 , \3478 , \3479 , \3480 , \3481 , \3482 , \3483 , \3484 , \3485 ,         \3486 , \3487 , \3488 , \3489 , \3490 , \3491 , \3492 , \3493 , \3494 , \3495 ,         \3496 , \3497 , \3498 , \3499 , \3500 , \3501 , \3502 , \3503 , \3504 , \3505 ,         \3506 , \3507 , \3508 , \3509 , \3510 , \3511 , \3512 , \3513 , \3514 , \3515 ,         \3516 , \3517 , \3518 , \3519 , \3520 , \3521 , \3522 , \3523 , \3524 , \3525 ,         \3526 , \3527 , \3528 , \3529 , \3530 , \3531 , \3532 , \3533 , \3534 , \3535 ,         \3536 , \3537 , \3538 , \3539 , \3540 , \3541 , \3542 , \3543 , \3544 , \3545 ,         \3546 , \3547 , \3548 , \3549 , \3550 , \3551 , \3552 , \3553 , \3554 , \3555 ,         \3556 , \3557 , \3558 , \3559 , \3560 , \3561 , \3562 , \3563 , \3564 , \3565 ,         \3566 , \3567 , \3568 , \3569 , \3570 , \3571 , \3572 , \3573 , \3574 , \3575 ,         \3576 , \3577 , \3578 , \3579 , \3580 , \3581 , \3582 , \3583 , \3584 , \3585 ,         \3586 , \3587 , \3588 , \3589 , \3590 , \3591 , \3592 , \3593 , \3594 , \3595 ,         \3596 , \3597 , \3598 , \3599 , \3600 , \3601 , \3602 , \3603 , \3604 , \3605 ,         \3606 , \3607 , \3608 , \3609 , \3610 , \3611 , \3612 , \3613 , \3614 , \3615 ,         \3616 , \3617 , \3618 , \3619 , \3620 , \3621 , \3622 , \3623 , \3624 , \3625 ,         \3626 , \3627 , \3628 , \3629 , \3630 , \3631 , \3632 , \3633 , \3634 , \3635 ,         \3636 , \3637 , \3638 , \3639 , \3640 , \3641 , \3642 , \3643 , \3644 , \3645 ,         \3646 , \3647 , \3648 , \3649 , \3650 , \3651 , \3652 , \3653 , \3654 , \3655 ,         \3656 , \3657 , \3658 , \3659 , \3660 , \3661 , \3662 , \3663 , \3664 , \3665 ,         \3666 , \3667 , \3668 , \3669 , \3670 , \3671 , \3672 , \3673 , \3674 , \3675 ,         \3676 , \3677 , \3678 , \3679 , \3680 , \3681 , \3682 , \3683 , \3684 , \3685 ,         \3686 , \3687 , \3688 , \3689 , \3690 , \3691 , \3692 , \3693 , \3694 , \3695 ,         \3696 , \3697 , \3698 , \3699 , \3700 , \3701 , \3702 , \3703 , \3704 , \3705 ,         \3706 , \3707 , \3708 , \3709 , \3710 , \3711 , \3712 , \3713 , \3714 , \3715 ,         \3716 , \3717 , \3718 , \3719 , \3720 , \3721 , \3722 , \3723 , \3724 , \3725 ,         \3726 , \3727 , \3728 , \3729 , \3730 , \3731 , \3732 , \3733 , \3734 , \3735 ,         \3736 , \3737 , \3738 , \3739 , \3740 , \3741 , \3742 , \3743 , \3744 , \3745 ,         \3746 , \3747 , \3748 , \3749 , \3750 , \3751 , \3752 , \3753 , \3754 , \3755 ,         \3756 , \3757 , \3758 , \3759 , \3760 , \3761 , \3762 , \3763 , \3764 , \3765 ,         \3766 , \3767 , \3768 , \3769 , \3770 , \3771 , \3772 , \3773 , \3774 , \3775 ,         \3776 , \3777 , \3778 , \3779 , \3780 , \3781 , \3782 , \3783 , \3784 , \3785 ,         \3786 , \3787 , \3788 , \3789 , \3790 , \3791 , \3792 , \3793 , \3794 , \3795 ,         \3796 , \3797 , \3798 , \3799 , \3800 , \3801 , \3802 , \3803 , \3804 , \3805 ,         \3806 , \3807 , \3808 , \3809 , \3810 , \3811 , \3812 , \3813 , \3814 , \3815 ,         \3816 , \3817 , \3818 , \3819 , \3820 , \3821 , \3822 , \3823 , \3824 , \3825 ,         \3826 , \3827 , \3828 , \3829 , \3830 , \3831 , \3832 , \3833 , \3834 , \3835 ,         \3836 , \3837 , \3838 , \3839 , \3840 , \3841 , \3842 , \3843 , \3844 , \3845 ,         \3846 , \3847 , \3848 , \3849 , \3850 , \3851 , \3852 , \3853 , \3854 , \3855 ,         \3856 , \3857 , \3858 , \3859 , \3860 , \3861 , \3862 , \3863 , \3864 , \3865 ,         \3866 , \3867 , \3868 , \3869 , \3870 , \3871 , \3872 , \3873 , \3874 , \3875 ,         \3876 , \3877 , \3878 , \3879 , \3880 , \3881 , \3882 , \3883 , \3884 , \3885 ,         \3886 , \3887 , \3888 , \3889 , \3890 , \3891 , \3892 , \3893 , \3894 , \3895 ,         \3896 , \3897 , \3898 , \3899 , \3900 , \3901 , \3902 , \3903 , \3904 , \3905 ,         \3906 , \3907 , \3908 , \3909 , \3910 , \3911 , \3912 , \3913 , \3914 , \3915 ,         \3916 , \3917 , \3918 , \3919 , \3920 , \3921 , \3922 , \3923 , \3924 , \3925 ,         \3926 , \3927 , \3928 , \3929 , \3930 , \3931 , \3932 , \3933 , \3934 , \3935 ,         \3936 , \3937 , \3938 , \3939 , \3940 , \3941 , \3942 , \3943 , \3944 , \3945 ,         \3946 , \3947 , \3948 , \3949 , \3950 , \3951 , \3952 , \3953 , \3954 , \3955 ,         \3956 , \3957 , \3958 , \3959 , \3960 , \3961 , \3962 , \3963 , \3964 , \3965 ,         \3966 , \3967 , \3968 , \3969 , \3970 , \3971 , \3972 , \3973 , \3974 , \3975 ,         \3976 , \3977 , \3978 , \3979 , \3980 , \3981 , \3982 , \3983 , \3984 , \3985 ,         \3986 , \3987 , \3988 , \3989 , \3990 , \3991 , \3992 , \3993 , \3994 , \3995 ,         \3996 , \3997 , \3998 , \3999 , \4000 , \4001 , \4002 , \4003 , \4004 , \4005 ,         \4006 , \4007 , \4008 , \4009 , \4010 , \4011 , \4012 , \4013 , \4014 , \4015 ,         \4016 , \4017 , \4018 , \4019 , \4020 , \4021 , \4022 , \4023 , \4024 , \4025 ,         \4026 , \4027 , \4028 , \4029 , \4030 , \4031 , \4032 , \4033 , \4034 , \4035 ,         \4036 , \4037 , \4038 , \4039 , \4040 , \4041 , \4042 , \4043 , \4044 , \4045 ,         \4046 , \4047 , \4048 , \4049 , \4050 , \4051 , \4052 , \4053 , \4054 , \4055 ,         \4056 , \4057 , \4058 , \4059 , \4060 , \4061 , \4062 , \4063 , \4064 , \4065 ,         \4066 , \4067 , \4068 , \4069 , \4070 , \4071 , \4072 , \4073 , \4074 , \4075 ,         \4076 , \4077 , \4078 , \4079 , \4080 , \4081 , \4082 , \4083 , \4084 , \4085 ,         \4086 , \4087 , \4088 , \4089 , \4090 , \4091 , \4092 , \4093 , \4094 , \4095 ,         \4096 , \4097 , \4098 , \4099 , \4100 , \4101 , \4102 , \4103 , \4104 , \4105 ,         \4106 , \4107 , \4108 , \4109 , \4110 , \4111 , \4112 , \4113 , \4114 , \4115 ,         \4116 , \4117 , \4118 , \4119 , \4120 , \4121 , \4122 , \4123 , \4124 , \4125 ,         \4126 , \4127 , \4128 , \4129 , \4130 , \4131 , \4132 , \4133 , \4134 , \4135 ,         \4136 , \4137 , \4138 , \4139 , \4140 , \4141 , \4142 , \4143 , \4144 , \4145 ,         \4146 , \4147 , \4148 , \4149 , \4150 , \4151 , \4152 , \4153 , \4154 , \4155 ,         \4156 , \4157 , \4158 , \4159 , \4160 , \4161 , \4162 , \4163 , \4164 , \4165 ,         \4166 , \4167 , \4168 , \4169 , \4170 , \4171 , \4172 , \4173 , \4174 , \4175 ,         \4176 , \4177 , \4178 , \4179 , \4180 , \4181 , \4182 , \4183 , \4184 , \4185 ,         \4186 , \4187 , \4188 , \4189 , \4190 , \4191 , \4192 , \4193 , \4194 , \4195 ,         \4196 , \4197 , \4198 , \4199 , \4200 , \4201 , \4202 , \4203 , \4204 , \4205 ,         \4206 , \4207 , \4208 , \4209 , \4210 , \4211 , \4212 , \4213 , \4214 , \4215 ,         \4216 , \4217 , \4218 , \4219 , \4220 , \4221 , \4222 , \4223 , \4224 , \4225 ,         \4226 , \4227 , \4228 , \4229 , \4230 , \4231 , \4232 , \4233 , \4234 , \4235 ,         \4236 , \4237 , \4238 , \4239 , \4240 , \4241 , \4242 , \4243 , \4244 , \4245 ,         \4246 , \4247 , \4248 , \4249 , \4250 , \4251 , \4252 , \4253 , \4254 , \4255 ,         \4256 , \4257 , \4258 , \4259 , \4260 , \4261 , \4262 , \4263 , \4264 , \4265 ,         \4266 , \4267 , \4268 , \4269 , \4270 , \4271 , \4272 , \4273 , \4274 , \4275 ,         \4276 , \4277 , \4278 , \4279 , \4280 , \4281 , \4282 , \4283 , \4284 , \4285 ,         \4286 , \4287 , \4288 , \4289 , \4290 , \4291 , \4292 , \4293 , \4294 , \4295 ,         \4296 , \4297 , \4298 , \4299 , \4300 , \4301 , \4302 , \4303 , \4304 , \4305 ,         \4306 , \4307 , \4308 , \4309 , \4310 , \4311 , \4312 , \4313 , \4314 , \4315 ,         \4316 , \4317 , \4318 , \4319 , \4320 , \4321 , \4322 , \4323 , \4324 , \4325 ,         \4326 , \4327 , \4328 , \4329 , \4330 , \4331 , \4332 , \4333 , \4334 , \4335 ,         \4336 , \4337 , \4338 , \4339 , \4340 , \4341 , \4342 , \4343 , \4344 , \4345 ,         \4346 , \4347 , \4348 , \4349 , \4350 , \4351 , \4352 , \4353 , \4354 , \4355 ,         \4356 , \4357 , \4358 , \4359 , \4360 , \4361 , \4362 , \4363 , \4364 , \4365 ,         \4366 , \4367 , \4368 , \4369 , \4370 , \4371 , \4372 , \4373 , \4374 , \4375 ,         \4376 , \4377 , \4378 , \4379 , \4380 , \4381 , \4382 , \4383 , \4384 , \4385 ,         \4386 , \4387 , \4388 , \4389 , \4390 , \4391 , \4392 , \4393 , \4394 , \4395 ,         \4396 , \4397 , \4398 , \4399 , \4400 , \4401 , \4402 , \4403 , \4404 , \4405 ,         \4406 , \4407 , \4408 , \4409 , \4410 , \4411 , \4412 , \4413 , \4414 , \4415 ,         \4416 , \4417 , \4418 , \4419 , \4420 , \4421 , \4422 , \4423 , \4424 , \4425 ,         \4426 , \4427 , \4428 , \4429 , \4430 , \4431 , \4432 , \4433 , \4434 , \4435 ,         \4436 , \4437 , \4438 , \4439 , \4440 , \4441 , \4442 , \4443 , \4444 , \4445 ,         \4446 , \4447 , \4448 , \4449 , \4450 , \4451 , \4452 , \4453 , \4454 , \4455 ,         \4456 , \4457 , \4458 , \4459 , \4460 , \4461 , \4462 , \4463 , \4464 , \4465 ,         \4466 , \4467 , \4468_Z[31] , \4469 , \4470_Z[30] , \4471 , \4472_Z[29] , \4473 , \4474_Z[28] , \4475 ,         \4476_Z[27] , \4477 , \4478_Z[26] , \4479 , \4480_Z[25] , \4481 , \4482_Z[24] , \4483 , \4484_Z[23] , \4485 ,         \4486_Z[22] , \4487 , \4488_Z[21] , \4489 , \4490_Z[20] , \4491 , \4492_Z[19] , \4493 , \4494_Z[18] , \4495 ,         \4496_Z[17] , \4497 , \4498_Z[16] , \4499 , \4500_Z[15] , \4501 , \4502_Z[14] , \4503 , \4504_Z[13] , \4505 ,         \4506_Z[12] , \4507 , \4508_Z[11] , \4509 , \4510_Z[10] , \4511 , \4512_Z[9] , \4513 , \4514_Z[8] , \4515 ,         \4516_Z[7] , \4517 , \4518_Z[6] , \4519 , \4520_Z[5] , \4521 , \4522_Z[4] , \4523 , \4524_Z[3] , \4525 ,         \4526_Z[2] , \4527 , \4528_Z[1] , \4529 , \4530_Z[0] ;
mbuf \U$labaj470 ( \o[31] , \4468_Z[31] );
mbuf \U$labaj471 ( \o[30] , \4470_Z[30] );
mbuf \U$labaj472 ( \o[29] , \4472_Z[29] );
mbuf \U$labaj473 ( \o[28] , \4474_Z[28] );
mbuf \U$labaj474 ( \o[27] , \4476_Z[27] );
mbuf \U$labaj475 ( \o[26] , \4478_Z[26] );
mbuf \U$labaj476 ( \o[25] , \4480_Z[25] );
mbuf \U$labaj477 ( \o[24] , \4482_Z[24] );
mbuf \U$labaj478 ( \o[23] , \4484_Z[23] );
mbuf \U$labaj479 ( \o[22] , \4486_Z[22] );
mbuf \U$labaj480 ( \o[21] , \4488_Z[21] );
mbuf \U$labaj481 ( \o[20] , \4490_Z[20] );
mbuf \U$labaj482 ( \o[19] , \4492_Z[19] );
mbuf \U$labaj483 ( \o[18] , \4494_Z[18] );
mbuf \U$labaj484 ( \o[17] , \4496_Z[17] );
mbuf \U$labaj485 ( \o[16] , \4498_Z[16] );
mbuf \U$labaj486 ( \o[15] , \4500_Z[15] );
mbuf \U$labaj487 ( \o[14] , \4502_Z[14] );
mbuf \U$labaj488 ( \o[13] , \4504_Z[13] );
mbuf \U$labaj489 ( \o[12] , \4506_Z[12] );
mbuf \U$labaj490 ( \o[11] , \4508_Z[11] );
mbuf \U$labaj491 ( \o[10] , \4510_Z[10] );
mbuf \U$labaj492 ( \o[9] , \4512_Z[9] );
mbuf \U$labaj493 ( \o[8] , \4514_Z[8] );
mbuf \U$labaj494 ( \o[7] , \4516_Z[7] );
mbuf \U$labaj495 ( \o[6] , \4518_Z[6] );
mbuf \U$labaj496 ( \o[5] , \4520_Z[5] );
mbuf \U$labaj497 ( \o[4] , \4522_Z[4] );
mbuf \U$labaj498 ( \o[3] , \4524_Z[3] );
mbuf \U$labaj499 ( \o[2] , \4526_Z[2] );
mbuf \U$labaj500 ( \o[1] , \4528_Z[1] );
mbuf \U$labaj501 ( \o[0] , \4530_Z[0] );
mbuf \mul_6_11/A[0] ( \156_A[0] , \a[0] );
mbuf \mul_6_11/B[0] ( \157_B[0] , \b[0] );
mand \mul_6_11/U$1408 ( \158 , \156_A[0] , \157_B[0] );
mbuf \mul_6_11/Z[0] ( \159_Z[0] , \158 );
mnot \U$9 ( \160 , \159_Z[0] );
mbuf \mul_6_11/A[1] ( \161_A[1] , \a[1] );
mand \mul_6_11/U$1407 ( \162 , \161_A[1] , \157_B[0] );
mbuf \mul_6_11/B[1] ( \163_B[1] , \b[1] );
mand \mul_6_11/U$1392 ( \164 , \156_A[0] , \163_B[1] );
mxor \mul_6_11/U$1376 ( \165 , \162 , \164 );
mbuf \mul_6_11/Z[1] ( \166_Z[1] , \165 );
mbuf \mul_6_11/A[2] ( \167_A[2] , \a[2] );
mand \mul_6_11/U$1406 ( \168 , \167_A[2] , \157_B[0] );
mand \mul_6_11/U$1391 ( \169 , \161_A[1] , \163_B[1] );
mxor \mul_6_11/U$1374 ( \170 , \168 , \169 );
mand \mul_6_11/U$1375 ( \171 , \162 , \164 );
mxor \mul_6_11/U$1371 ( \172 , \170 , \171 );
mbuf \mul_6_11/B[2] ( \173_B[2] , \b[2] );
mand \mul_6_11/U$1302 ( \174 , \156_A[0] , \173_B[2] );
mxor \mul_6_11/U$1286 ( \175 , \172 , \174 );
mbuf \mul_6_11/Z[2] ( \176_Z[2] , \175 );
mbuf \mul_6_11/A[3] ( \177_A[3] , \a[3] );
mand \mul_6_11/U$1405 ( \178 , \177_A[3] , \157_B[0] );
mand \mul_6_11/U$1390 ( \179 , \167_A[2] , \163_B[1] );
mxor \mul_6_11/U$1369 ( \180 , \178 , \179 );
mand \mul_6_11/U$1373 ( \181 , \168 , \169 );
mand \mul_6_11/U$1372 ( \182 , \170 , \171 );
mor \mul_6_11/U$1370 ( \183 , \181 , \182 );
mxor \mul_6_11/U$1366 ( \184 , \180 , \183 );
mand \mul_6_11/U$1301 ( \185 , \161_A[1] , \173_B[2] );
mxor \mul_6_11/U$1284 ( \186 , \184 , \185 );
mand \mul_6_11/U$1285 ( \187 , \172 , \174 );
mxor \mul_6_11/U$1281 ( \188 , \186 , \187 );
mbuf \mul_6_11/B[3] ( \189_B[3] , \b[3] );
mand \mul_6_11/U$1209 ( \190 , \156_A[0] , \189_B[3] );
mxor \mul_6_11/U$1193 ( \191 , \188 , \190 );
mbuf \mul_6_11/Z[3] ( \192_Z[3] , \191 );
mbuf \mul_6_11/A[4] ( \193_A[4] , \a[4] );
mand \mul_6_11/U$1404 ( \194 , \193_A[4] , \157_B[0] );
mand \mul_6_11/U$1389 ( \195 , \177_A[3] , \163_B[1] );
mxor \mul_6_11/U$1364 ( \196 , \194 , \195 );
mand \mul_6_11/U$1368 ( \197 , \178 , \179 );
mand \mul_6_11/U$1367 ( \198 , \180 , \183 );
mor \mul_6_11/U$1365 ( \199 , \197 , \198 );
mxor \mul_6_11/U$1361 ( \200 , \196 , \199 );
mand \mul_6_11/U$1300 ( \201 , \167_A[2] , \173_B[2] );
mxor \mul_6_11/U$1279 ( \202 , \200 , \201 );
mand \mul_6_11/U$1283 ( \203 , \184 , \185 );
mand \mul_6_11/U$1282 ( \204 , \186 , \187 );
mor \mul_6_11/U$1280 ( \205 , \203 , \204 );
mxor \mul_6_11/U$1276 ( \206 , \202 , \205 );
mand \mul_6_11/U$1208 ( \207 , \161_A[1] , \189_B[3] );
mxor \mul_6_11/U$1191 ( \208 , \206 , \207 );
mand \mul_6_11/U$1192 ( \209 , \188 , \190 );
mxor \mul_6_11/U$1188 ( \210 , \208 , \209 );
mbuf \mul_6_11/B[4] ( \211_B[4] , \b[4] );
mand \mul_6_11/U$1116 ( \212 , \156_A[0] , \211_B[4] );
mxor \mul_6_11/U$1100 ( \213 , \210 , \212 );
mbuf \mul_6_11/Z[4] ( \214_Z[4] , \213 );
mbuf \mul_6_11/A[5] ( \215_A[5] , \a[5] );
mand \mul_6_11/U$1403 ( \216 , \215_A[5] , \157_B[0] );
mand \mul_6_11/U$1388 ( \217 , \193_A[4] , \163_B[1] );
mxor \mul_6_11/U$1359 ( \218 , \216 , \217 );
mand \mul_6_11/U$1363 ( \219 , \194 , \195 );
mand \mul_6_11/U$1362 ( \220 , \196 , \199 );
mor \mul_6_11/U$1360 ( \221 , \219 , \220 );
mxor \mul_6_11/U$1356 ( \222 , \218 , \221 );
mand \mul_6_11/U$1299 ( \223 , \177_A[3] , \173_B[2] );
mxor \mul_6_11/U$1274 ( \224 , \222 , \223 );
mand \mul_6_11/U$1278 ( \225 , \200 , \201 );
mand \mul_6_11/U$1277 ( \226 , \202 , \205 );
mor \mul_6_11/U$1275 ( \227 , \225 , \226 );
mxor \mul_6_11/U$1271 ( \228 , \224 , \227 );
mand \mul_6_11/U$1207 ( \229 , \167_A[2] , \189_B[3] );
mxor \mul_6_11/U$1186 ( \230 , \228 , \229 );
mand \mul_6_11/U$1190 ( \231 , \206 , \207 );
mand \mul_6_11/U$1189 ( \232 , \208 , \209 );
mor \mul_6_11/U$1187 ( \233 , \231 , \232 );
mxor \mul_6_11/U$1183 ( \234 , \230 , \233 );
mand \mul_6_11/U$1115 ( \235 , \161_A[1] , \211_B[4] );
mxor \mul_6_11/U$1098 ( \236 , \234 , \235 );
mand \mul_6_11/U$1099 ( \237 , \210 , \212 );
mxor \mul_6_11/U$1095 ( \238 , \236 , \237 );
mbuf \mul_6_11/B[5] ( \239_B[5] , \b[5] );
mand \mul_6_11/U$1023 ( \240 , \156_A[0] , \239_B[5] );
mxor \mul_6_11/U$1007 ( \241 , \238 , \240 );
mbuf \mul_6_11/Z[5] ( \242_Z[5] , \241 );
mbuf \mul_6_11/A[6] ( \243_A[6] , \a[6] );
mand \mul_6_11/U$1402 ( \244 , \243_A[6] , \157_B[0] );
mand \mul_6_11/U$1387 ( \245 , \215_A[5] , \163_B[1] );
mxor \mul_6_11/U$1354 ( \246 , \244 , \245 );
mand \mul_6_11/U$1358 ( \247 , \216 , \217 );
mand \mul_6_11/U$1357 ( \248 , \218 , \221 );
mor \mul_6_11/U$1355 ( \249 , \247 , \248 );
mxor \mul_6_11/U$1351 ( \250 , \246 , \249 );
mand \mul_6_11/U$1298 ( \251 , \193_A[4] , \173_B[2] );
mxor \mul_6_11/U$1269 ( \252 , \250 , \251 );
mand \mul_6_11/U$1273 ( \253 , \222 , \223 );
mand \mul_6_11/U$1272 ( \254 , \224 , \227 );
mor \mul_6_11/U$1270 ( \255 , \253 , \254 );
mxor \mul_6_11/U$1266 ( \256 , \252 , \255 );
mand \mul_6_11/U$1206 ( \257 , \177_A[3] , \189_B[3] );
mxor \mul_6_11/U$1181 ( \258 , \256 , \257 );
mand \mul_6_11/U$1185 ( \259 , \228 , \229 );
mand \mul_6_11/U$1184 ( \260 , \230 , \233 );
mor \mul_6_11/U$1182 ( \261 , \259 , \260 );
mxor \mul_6_11/U$1178 ( \262 , \258 , \261 );
mand \mul_6_11/U$1114 ( \263 , \167_A[2] , \211_B[4] );
mxor \mul_6_11/U$1093 ( \264 , \262 , \263 );
mand \mul_6_11/U$1097 ( \265 , \234 , \235 );
mand \mul_6_11/U$1096 ( \266 , \236 , \237 );
mor \mul_6_11/U$1094 ( \267 , \265 , \266 );
mxor \mul_6_11/U$1090 ( \268 , \264 , \267 );
mand \mul_6_11/U$1022 ( \269 , \161_A[1] , \239_B[5] );
mxor \mul_6_11/U$1005 ( \270 , \268 , \269 );
mand \mul_6_11/U$1006 ( \271 , \238 , \240 );
mxor \mul_6_11/U$1002 ( \272 , \270 , \271 );
mbuf \mul_6_11/B[6] ( \273_B[6] , \b[6] );
mand \mul_6_11/U$930 ( \274 , \156_A[0] , \273_B[6] );
mxor \mul_6_11/U$914 ( \275 , \272 , \274 );
mbuf \mul_6_11/Z[6] ( \276_Z[6] , \275 );
mbuf \mul_6_11/A[7] ( \277_A[7] , \a[7] );
mand \mul_6_11/U$1401 ( \278 , \277_A[7] , \157_B[0] );
mand \mul_6_11/U$1386 ( \279 , \243_A[6] , \163_B[1] );
mxor \mul_6_11/U$1349 ( \280 , \278 , \279 );
mand \mul_6_11/U$1353 ( \281 , \244 , \245 );
mand \mul_6_11/U$1352 ( \282 , \246 , \249 );
mor \mul_6_11/U$1350 ( \283 , \281 , \282 );
mxor \mul_6_11/U$1346 ( \284 , \280 , \283 );
mand \mul_6_11/U$1297 ( \285 , \215_A[5] , \173_B[2] );
mxor \mul_6_11/U$1264 ( \286 , \284 , \285 );
mand \mul_6_11/U$1268 ( \287 , \250 , \251 );
mand \mul_6_11/U$1267 ( \288 , \252 , \255 );
mor \mul_6_11/U$1265 ( \289 , \287 , \288 );
mxor \mul_6_11/U$1261 ( \290 , \286 , \289 );
mand \mul_6_11/U$1205 ( \291 , \193_A[4] , \189_B[3] );
mxor \mul_6_11/U$1176 ( \292 , \290 , \291 );
mand \mul_6_11/U$1180 ( \293 , \256 , \257 );
mand \mul_6_11/U$1179 ( \294 , \258 , \261 );
mor \mul_6_11/U$1177 ( \295 , \293 , \294 );
mxor \mul_6_11/U$1173 ( \296 , \292 , \295 );
mand \mul_6_11/U$1113 ( \297 , \177_A[3] , \211_B[4] );
mxor \mul_6_11/U$1088 ( \298 , \296 , \297 );
mand \mul_6_11/U$1092 ( \299 , \262 , \263 );
mand \mul_6_11/U$1091 ( \300 , \264 , \267 );
mor \mul_6_11/U$1089 ( \301 , \299 , \300 );
mxor \mul_6_11/U$1085 ( \302 , \298 , \301 );
mand \mul_6_11/U$1021 ( \303 , \167_A[2] , \239_B[5] );
mxor \mul_6_11/U$1000 ( \304 , \302 , \303 );
mand \mul_6_11/U$1004 ( \305 , \268 , \269 );
mand \mul_6_11/U$1003 ( \306 , \270 , \271 );
mor \mul_6_11/U$1001 ( \307 , \305 , \306 );
mxor \mul_6_11/U$997 ( \308 , \304 , \307 );
mand \mul_6_11/U$929 ( \309 , \161_A[1] , \273_B[6] );
mxor \mul_6_11/U$912 ( \310 , \308 , \309 );
mand \mul_6_11/U$913 ( \311 , \272 , \274 );
mxor \mul_6_11/U$909 ( \312 , \310 , \311 );
mbuf \mul_6_11/B[7] ( \313_B[7] , \b[7] );
mand \mul_6_11/U$837 ( \314 , \156_A[0] , \313_B[7] );
mxor \mul_6_11/U$821 ( \315 , \312 , \314 );
mbuf \mul_6_11/Z[7] ( \316_Z[7] , \315 );
mbuf \mul_6_11/A[8] ( \317_A[8] , \a[8] );
mand \mul_6_11/U$1400 ( \318 , \317_A[8] , \157_B[0] );
mand \mul_6_11/U$1385 ( \319 , \277_A[7] , \163_B[1] );
mxor \mul_6_11/U$1344 ( \320 , \318 , \319 );
mand \mul_6_11/U$1348 ( \321 , \278 , \279 );
mand \mul_6_11/U$1347 ( \322 , \280 , \283 );
mor \mul_6_11/U$1345 ( \323 , \321 , \322 );
mxor \mul_6_11/U$1341 ( \324 , \320 , \323 );
mand \mul_6_11/U$1296 ( \325 , \243_A[6] , \173_B[2] );
mxor \mul_6_11/U$1259 ( \326 , \324 , \325 );
mand \mul_6_11/U$1263 ( \327 , \284 , \285 );
mand \mul_6_11/U$1262 ( \328 , \286 , \289 );
mor \mul_6_11/U$1260 ( \329 , \327 , \328 );
mxor \mul_6_11/U$1256 ( \330 , \326 , \329 );
mand \mul_6_11/U$1204 ( \331 , \215_A[5] , \189_B[3] );
mxor \mul_6_11/U$1171 ( \332 , \330 , \331 );
mand \mul_6_11/U$1175 ( \333 , \290 , \291 );
mand \mul_6_11/U$1174 ( \334 , \292 , \295 );
mor \mul_6_11/U$1172 ( \335 , \333 , \334 );
mxor \mul_6_11/U$1168 ( \336 , \332 , \335 );
mand \mul_6_11/U$1112 ( \337 , \193_A[4] , \211_B[4] );
mxor \mul_6_11/U$1083 ( \338 , \336 , \337 );
mand \mul_6_11/U$1087 ( \339 , \296 , \297 );
mand \mul_6_11/U$1086 ( \340 , \298 , \301 );
mor \mul_6_11/U$1084 ( \341 , \339 , \340 );
mxor \mul_6_11/U$1080 ( \342 , \338 , \341 );
mand \mul_6_11/U$1020 ( \343 , \177_A[3] , \239_B[5] );
mxor \mul_6_11/U$995 ( \344 , \342 , \343 );
mand \mul_6_11/U$999 ( \345 , \302 , \303 );
mand \mul_6_11/U$998 ( \346 , \304 , \307 );
mor \mul_6_11/U$996 ( \347 , \345 , \346 );
mxor \mul_6_11/U$992 ( \348 , \344 , \347 );
mand \mul_6_11/U$928 ( \349 , \167_A[2] , \273_B[6] );
mxor \mul_6_11/U$907 ( \350 , \348 , \349 );
mand \mul_6_11/U$911 ( \351 , \308 , \309 );
mand \mul_6_11/U$910 ( \352 , \310 , \311 );
mor \mul_6_11/U$908 ( \353 , \351 , \352 );
mxor \mul_6_11/U$904 ( \354 , \350 , \353 );
mand \mul_6_11/U$836 ( \355 , \161_A[1] , \313_B[7] );
mxor \mul_6_11/U$819 ( \356 , \354 , \355 );
mand \mul_6_11/U$820 ( \357 , \312 , \314 );
mxor \mul_6_11/U$816 ( \358 , \356 , \357 );
mbuf \mul_6_11/B[8] ( \359_B[8] , \b[8] );
mand \mul_6_11/U$744 ( \360 , \156_A[0] , \359_B[8] );
mxor \mul_6_11/U$728 ( \361 , \358 , \360 );
mbuf \mul_6_11/Z[8] ( \362_Z[8] , \361 );
mbuf \mul_6_11/A[9] ( \363_A[9] , \a[9] );
mand \mul_6_11/U$1399 ( \364 , \363_A[9] , \157_B[0] );
mand \mul_6_11/U$1384 ( \365 , \317_A[8] , \163_B[1] );
mxor \mul_6_11/U$1339 ( \366 , \364 , \365 );
mand \mul_6_11/U$1343 ( \367 , \318 , \319 );
mand \mul_6_11/U$1342 ( \368 , \320 , \323 );
mor \mul_6_11/U$1340 ( \369 , \367 , \368 );
mxor \mul_6_11/U$1336 ( \370 , \366 , \369 );
mand \mul_6_11/U$1295 ( \371 , \277_A[7] , \173_B[2] );
mxor \mul_6_11/U$1254 ( \372 , \370 , \371 );
mand \mul_6_11/U$1258 ( \373 , \324 , \325 );
mand \mul_6_11/U$1257 ( \374 , \326 , \329 );
mor \mul_6_11/U$1255 ( \375 , \373 , \374 );
mxor \mul_6_11/U$1251 ( \376 , \372 , \375 );
mand \mul_6_11/U$1203 ( \377 , \243_A[6] , \189_B[3] );
mxor \mul_6_11/U$1166 ( \378 , \376 , \377 );
mand \mul_6_11/U$1170 ( \379 , \330 , \331 );
mand \mul_6_11/U$1169 ( \380 , \332 , \335 );
mor \mul_6_11/U$1167 ( \381 , \379 , \380 );
mxor \mul_6_11/U$1163 ( \382 , \378 , \381 );
mand \mul_6_11/U$1111 ( \383 , \215_A[5] , \211_B[4] );
mxor \mul_6_11/U$1078 ( \384 , \382 , \383 );
mand \mul_6_11/U$1082 ( \385 , \336 , \337 );
mand \mul_6_11/U$1081 ( \386 , \338 , \341 );
mor \mul_6_11/U$1079 ( \387 , \385 , \386 );
mxor \mul_6_11/U$1075 ( \388 , \384 , \387 );
mand \mul_6_11/U$1019 ( \389 , \193_A[4] , \239_B[5] );
mxor \mul_6_11/U$990 ( \390 , \388 , \389 );
mand \mul_6_11/U$994 ( \391 , \342 , \343 );
mand \mul_6_11/U$993 ( \392 , \344 , \347 );
mor \mul_6_11/U$991 ( \393 , \391 , \392 );
mxor \mul_6_11/U$987 ( \394 , \390 , \393 );
mand \mul_6_11/U$927 ( \395 , \177_A[3] , \273_B[6] );
mxor \mul_6_11/U$902 ( \396 , \394 , \395 );
mand \mul_6_11/U$906 ( \397 , \348 , \349 );
mand \mul_6_11/U$905 ( \398 , \350 , \353 );
mor \mul_6_11/U$903 ( \399 , \397 , \398 );
mxor \mul_6_11/U$899 ( \400 , \396 , \399 );
mand \mul_6_11/U$835 ( \401 , \167_A[2] , \313_B[7] );
mxor \mul_6_11/U$814 ( \402 , \400 , \401 );
mand \mul_6_11/U$818 ( \403 , \354 , \355 );
mand \mul_6_11/U$817 ( \404 , \356 , \357 );
mor \mul_6_11/U$815 ( \405 , \403 , \404 );
mxor \mul_6_11/U$811 ( \406 , \402 , \405 );
mand \mul_6_11/U$743 ( \407 , \161_A[1] , \359_B[8] );
mxor \mul_6_11/U$726 ( \408 , \406 , \407 );
mand \mul_6_11/U$727 ( \409 , \358 , \360 );
mxor \mul_6_11/U$723 ( \410 , \408 , \409 );
mbuf \mul_6_11/B[9] ( \411_B[9] , \b[9] );
mand \mul_6_11/U$651 ( \412 , \156_A[0] , \411_B[9] );
mxor \mul_6_11/U$635 ( \413 , \410 , \412 );
mbuf \mul_6_11/Z[9] ( \414_Z[9] , \413 );
mbuf \mul_6_11/A[10] ( \415_A[10] , \a[10] );
mand \mul_6_11/U$1398 ( \416 , \415_A[10] , \157_B[0] );
mand \mul_6_11/U$1383 ( \417 , \363_A[9] , \163_B[1] );
mxor \mul_6_11/U$1334 ( \418 , \416 , \417 );
mand \mul_6_11/U$1338 ( \419 , \364 , \365 );
mand \mul_6_11/U$1337 ( \420 , \366 , \369 );
mor \mul_6_11/U$1335 ( \421 , \419 , \420 );
mxor \mul_6_11/U$1331 ( \422 , \418 , \421 );
mand \mul_6_11/U$1294 ( \423 , \317_A[8] , \173_B[2] );
mxor \mul_6_11/U$1249 ( \424 , \422 , \423 );
mand \mul_6_11/U$1253 ( \425 , \370 , \371 );
mand \mul_6_11/U$1252 ( \426 , \372 , \375 );
mor \mul_6_11/U$1250 ( \427 , \425 , \426 );
mxor \mul_6_11/U$1246 ( \428 , \424 , \427 );
mand \mul_6_11/U$1202 ( \429 , \277_A[7] , \189_B[3] );
mxor \mul_6_11/U$1161 ( \430 , \428 , \429 );
mand \mul_6_11/U$1165 ( \431 , \376 , \377 );
mand \mul_6_11/U$1164 ( \432 , \378 , \381 );
mor \mul_6_11/U$1162 ( \433 , \431 , \432 );
mxor \mul_6_11/U$1158 ( \434 , \430 , \433 );
mand \mul_6_11/U$1110 ( \435 , \243_A[6] , \211_B[4] );
mxor \mul_6_11/U$1073 ( \436 , \434 , \435 );
mand \mul_6_11/U$1077 ( \437 , \382 , \383 );
mand \mul_6_11/U$1076 ( \438 , \384 , \387 );
mor \mul_6_11/U$1074 ( \439 , \437 , \438 );
mxor \mul_6_11/U$1070 ( \440 , \436 , \439 );
mand \mul_6_11/U$1018 ( \441 , \215_A[5] , \239_B[5] );
mxor \mul_6_11/U$985 ( \442 , \440 , \441 );
mand \mul_6_11/U$989 ( \443 , \388 , \389 );
mand \mul_6_11/U$988 ( \444 , \390 , \393 );
mor \mul_6_11/U$986 ( \445 , \443 , \444 );
mxor \mul_6_11/U$982 ( \446 , \442 , \445 );
mand \mul_6_11/U$926 ( \447 , \193_A[4] , \273_B[6] );
mxor \mul_6_11/U$897 ( \448 , \446 , \447 );
mand \mul_6_11/U$901 ( \449 , \394 , \395 );
mand \mul_6_11/U$900 ( \450 , \396 , \399 );
mor \mul_6_11/U$898 ( \451 , \449 , \450 );
mxor \mul_6_11/U$894 ( \452 , \448 , \451 );
mand \mul_6_11/U$834 ( \453 , \177_A[3] , \313_B[7] );
mxor \mul_6_11/U$809 ( \454 , \452 , \453 );
mand \mul_6_11/U$813 ( \455 , \400 , \401 );
mand \mul_6_11/U$812 ( \456 , \402 , \405 );
mor \mul_6_11/U$810 ( \457 , \455 , \456 );
mxor \mul_6_11/U$806 ( \458 , \454 , \457 );
mand \mul_6_11/U$742 ( \459 , \167_A[2] , \359_B[8] );
mxor \mul_6_11/U$721 ( \460 , \458 , \459 );
mand \mul_6_11/U$725 ( \461 , \406 , \407 );
mand \mul_6_11/U$724 ( \462 , \408 , \409 );
mor \mul_6_11/U$722 ( \463 , \461 , \462 );
mxor \mul_6_11/U$718 ( \464 , \460 , \463 );
mand \mul_6_11/U$650 ( \465 , \161_A[1] , \411_B[9] );
mxor \mul_6_11/U$633 ( \466 , \464 , \465 );
mand \mul_6_11/U$634 ( \467 , \410 , \412 );
mxor \mul_6_11/U$630 ( \468 , \466 , \467 );
mbuf \mul_6_11/B[10] ( \469_B[10] , \b[10] );
mand \mul_6_11/U$558 ( \470 , \156_A[0] , \469_B[10] );
mxor \mul_6_11/U$542 ( \471 , \468 , \470 );
mbuf \mul_6_11/Z[10] ( \472_Z[10] , \471 );
mbuf \mul_6_11/A[11] ( \473_A[11] , \a[11] );
mand \mul_6_11/U$1397 ( \474 , \473_A[11] , \157_B[0] );
mand \mul_6_11/U$1382 ( \475 , \415_A[10] , \163_B[1] );
mxor \mul_6_11/U$1329 ( \476 , \474 , \475 );
mand \mul_6_11/U$1333 ( \477 , \416 , \417 );
mand \mul_6_11/U$1332 ( \478 , \418 , \421 );
mor \mul_6_11/U$1330 ( \479 , \477 , \478 );
mxor \mul_6_11/U$1326 ( \480 , \476 , \479 );
mand \mul_6_11/U$1293 ( \481 , \363_A[9] , \173_B[2] );
mxor \mul_6_11/U$1244 ( \482 , \480 , \481 );
mand \mul_6_11/U$1248 ( \483 , \422 , \423 );
mand \mul_6_11/U$1247 ( \484 , \424 , \427 );
mor \mul_6_11/U$1245 ( \485 , \483 , \484 );
mxor \mul_6_11/U$1241 ( \486 , \482 , \485 );
mand \mul_6_11/U$1201 ( \487 , \317_A[8] , \189_B[3] );
mxor \mul_6_11/U$1156 ( \488 , \486 , \487 );
mand \mul_6_11/U$1160 ( \489 , \428 , \429 );
mand \mul_6_11/U$1159 ( \490 , \430 , \433 );
mor \mul_6_11/U$1157 ( \491 , \489 , \490 );
mxor \mul_6_11/U$1153 ( \492 , \488 , \491 );
mand \mul_6_11/U$1109 ( \493 , \277_A[7] , \211_B[4] );
mxor \mul_6_11/U$1068 ( \494 , \492 , \493 );
mand \mul_6_11/U$1072 ( \495 , \434 , \435 );
mand \mul_6_11/U$1071 ( \496 , \436 , \439 );
mor \mul_6_11/U$1069 ( \497 , \495 , \496 );
mxor \mul_6_11/U$1065 ( \498 , \494 , \497 );
mand \mul_6_11/U$1017 ( \499 , \243_A[6] , \239_B[5] );
mxor \mul_6_11/U$980 ( \500 , \498 , \499 );
mand \mul_6_11/U$984 ( \501 , \440 , \441 );
mand \mul_6_11/U$983 ( \502 , \442 , \445 );
mor \mul_6_11/U$981 ( \503 , \501 , \502 );
mxor \mul_6_11/U$977 ( \504 , \500 , \503 );
mand \mul_6_11/U$925 ( \505 , \215_A[5] , \273_B[6] );
mxor \mul_6_11/U$892 ( \506 , \504 , \505 );
mand \mul_6_11/U$896 ( \507 , \446 , \447 );
mand \mul_6_11/U$895 ( \508 , \448 , \451 );
mor \mul_6_11/U$893 ( \509 , \507 , \508 );
mxor \mul_6_11/U$889 ( \510 , \506 , \509 );
mand \mul_6_11/U$833 ( \511 , \193_A[4] , \313_B[7] );
mxor \mul_6_11/U$804 ( \512 , \510 , \511 );
mand \mul_6_11/U$808 ( \513 , \452 , \453 );
mand \mul_6_11/U$807 ( \514 , \454 , \457 );
mor \mul_6_11/U$805 ( \515 , \513 , \514 );
mxor \mul_6_11/U$801 ( \516 , \512 , \515 );
mand \mul_6_11/U$741 ( \517 , \177_A[3] , \359_B[8] );
mxor \mul_6_11/U$716 ( \518 , \516 , \517 );
mand \mul_6_11/U$720 ( \519 , \458 , \459 );
mand \mul_6_11/U$719 ( \520 , \460 , \463 );
mor \mul_6_11/U$717 ( \521 , \519 , \520 );
mxor \mul_6_11/U$713 ( \522 , \518 , \521 );
mand \mul_6_11/U$649 ( \523 , \167_A[2] , \411_B[9] );
mxor \mul_6_11/U$628 ( \524 , \522 , \523 );
mand \mul_6_11/U$632 ( \525 , \464 , \465 );
mand \mul_6_11/U$631 ( \526 , \466 , \467 );
mor \mul_6_11/U$629 ( \527 , \525 , \526 );
mxor \mul_6_11/U$625 ( \528 , \524 , \527 );
mand \mul_6_11/U$557 ( \529 , \161_A[1] , \469_B[10] );
mxor \mul_6_11/U$540 ( \530 , \528 , \529 );
mand \mul_6_11/U$541 ( \531 , \468 , \470 );
mxor \mul_6_11/U$537 ( \532 , \530 , \531 );
mbuf \mul_6_11/B[11] ( \533_B[11] , \b[11] );
mand \mul_6_11/U$465 ( \534 , \156_A[0] , \533_B[11] );
mxor \mul_6_11/U$449 ( \535 , \532 , \534 );
mbuf \mul_6_11/Z[11] ( \536_Z[11] , \535 );
mbuf \mul_6_11/A[12] ( \537_A[12] , \a[12] );
mand \mul_6_11/U$1396 ( \538 , \537_A[12] , \157_B[0] );
mand \mul_6_11/U$1381 ( \539 , \473_A[11] , \163_B[1] );
mxor \mul_6_11/U$1324 ( \540 , \538 , \539 );
mand \mul_6_11/U$1328 ( \541 , \474 , \475 );
mand \mul_6_11/U$1327 ( \542 , \476 , \479 );
mor \mul_6_11/U$1325 ( \543 , \541 , \542 );
mxor \mul_6_11/U$1321 ( \544 , \540 , \543 );
mand \mul_6_11/U$1292 ( \545 , \415_A[10] , \173_B[2] );
mxor \mul_6_11/U$1239 ( \546 , \544 , \545 );
mand \mul_6_11/U$1243 ( \547 , \480 , \481 );
mand \mul_6_11/U$1242 ( \548 , \482 , \485 );
mor \mul_6_11/U$1240 ( \549 , \547 , \548 );
mxor \mul_6_11/U$1236 ( \550 , \546 , \549 );
mand \mul_6_11/U$1200 ( \551 , \363_A[9] , \189_B[3] );
mxor \mul_6_11/U$1151 ( \552 , \550 , \551 );
mand \mul_6_11/U$1155 ( \553 , \486 , \487 );
mand \mul_6_11/U$1154 ( \554 , \488 , \491 );
mor \mul_6_11/U$1152 ( \555 , \553 , \554 );
mxor \mul_6_11/U$1148 ( \556 , \552 , \555 );
mand \mul_6_11/U$1108 ( \557 , \317_A[8] , \211_B[4] );
mxor \mul_6_11/U$1063 ( \558 , \556 , \557 );
mand \mul_6_11/U$1067 ( \559 , \492 , \493 );
mand \mul_6_11/U$1066 ( \560 , \494 , \497 );
mor \mul_6_11/U$1064 ( \561 , \559 , \560 );
mxor \mul_6_11/U$1060 ( \562 , \558 , \561 );
mand \mul_6_11/U$1016 ( \563 , \277_A[7] , \239_B[5] );
mxor \mul_6_11/U$975 ( \564 , \562 , \563 );
mand \mul_6_11/U$979 ( \565 , \498 , \499 );
mand \mul_6_11/U$978 ( \566 , \500 , \503 );
mor \mul_6_11/U$976 ( \567 , \565 , \566 );
mxor \mul_6_11/U$972 ( \568 , \564 , \567 );
mand \mul_6_11/U$924 ( \569 , \243_A[6] , \273_B[6] );
mxor \mul_6_11/U$887 ( \570 , \568 , \569 );
mand \mul_6_11/U$891 ( \571 , \504 , \505 );
mand \mul_6_11/U$890 ( \572 , \506 , \509 );
mor \mul_6_11/U$888 ( \573 , \571 , \572 );
mxor \mul_6_11/U$884 ( \574 , \570 , \573 );
mand \mul_6_11/U$832 ( \575 , \215_A[5] , \313_B[7] );
mxor \mul_6_11/U$799 ( \576 , \574 , \575 );
mand \mul_6_11/U$803 ( \577 , \510 , \511 );
mand \mul_6_11/U$802 ( \578 , \512 , \515 );
mor \mul_6_11/U$800 ( \579 , \577 , \578 );
mxor \mul_6_11/U$796 ( \580 , \576 , \579 );
mand \mul_6_11/U$740 ( \581 , \193_A[4] , \359_B[8] );
mxor \mul_6_11/U$711 ( \582 , \580 , \581 );
mand \mul_6_11/U$715 ( \583 , \516 , \517 );
mand \mul_6_11/U$714 ( \584 , \518 , \521 );
mor \mul_6_11/U$712 ( \585 , \583 , \584 );
mxor \mul_6_11/U$708 ( \586 , \582 , \585 );
mand \mul_6_11/U$648 ( \587 , \177_A[3] , \411_B[9] );
mxor \mul_6_11/U$623 ( \588 , \586 , \587 );
mand \mul_6_11/U$627 ( \589 , \522 , \523 );
mand \mul_6_11/U$626 ( \590 , \524 , \527 );
mor \mul_6_11/U$624 ( \591 , \589 , \590 );
mxor \mul_6_11/U$620 ( \592 , \588 , \591 );
mand \mul_6_11/U$556 ( \593 , \167_A[2] , \469_B[10] );
mxor \mul_6_11/U$535 ( \594 , \592 , \593 );
mand \mul_6_11/U$539 ( \595 , \528 , \529 );
mand \mul_6_11/U$538 ( \596 , \530 , \531 );
mor \mul_6_11/U$536 ( \597 , \595 , \596 );
mxor \mul_6_11/U$532 ( \598 , \594 , \597 );
mand \mul_6_11/U$464 ( \599 , \161_A[1] , \533_B[11] );
mxor \mul_6_11/U$447 ( \600 , \598 , \599 );
mand \mul_6_11/U$448 ( \601 , \532 , \534 );
mxor \mul_6_11/U$444 ( \602 , \600 , \601 );
mbuf \mul_6_11/B[12] ( \603_B[12] , \b[12] );
mand \mul_6_11/U$372 ( \604 , \156_A[0] , \603_B[12] );
mxor \mul_6_11/U$356 ( \605 , \602 , \604 );
mbuf \mul_6_11/Z[12] ( \606_Z[12] , \605 );
mbuf \mul_6_11/A[13] ( \607_A[13] , \a[13] );
mand \mul_6_11/U$1395 ( \608 , \607_A[13] , \157_B[0] );
mand \mul_6_11/U$1380 ( \609 , \537_A[12] , \163_B[1] );
mxor \mul_6_11/U$1319 ( \610 , \608 , \609 );
mand \mul_6_11/U$1323 ( \611 , \538 , \539 );
mand \mul_6_11/U$1322 ( \612 , \540 , \543 );
mor \mul_6_11/U$1320 ( \613 , \611 , \612 );
mxor \mul_6_11/U$1316 ( \614 , \610 , \613 );
mand \mul_6_11/U$1291 ( \615 , \473_A[11] , \173_B[2] );
mxor \mul_6_11/U$1234 ( \616 , \614 , \615 );
mand \mul_6_11/U$1238 ( \617 , \544 , \545 );
mand \mul_6_11/U$1237 ( \618 , \546 , \549 );
mor \mul_6_11/U$1235 ( \619 , \617 , \618 );
mxor \mul_6_11/U$1231 ( \620 , \616 , \619 );
mand \mul_6_11/U$1199 ( \621 , \415_A[10] , \189_B[3] );
mxor \mul_6_11/U$1146 ( \622 , \620 , \621 );
mand \mul_6_11/U$1150 ( \623 , \550 , \551 );
mand \mul_6_11/U$1149 ( \624 , \552 , \555 );
mor \mul_6_11/U$1147 ( \625 , \623 , \624 );
mxor \mul_6_11/U$1143 ( \626 , \622 , \625 );
mand \mul_6_11/U$1107 ( \627 , \363_A[9] , \211_B[4] );
mxor \mul_6_11/U$1058 ( \628 , \626 , \627 );
mand \mul_6_11/U$1062 ( \629 , \556 , \557 );
mand \mul_6_11/U$1061 ( \630 , \558 , \561 );
mor \mul_6_11/U$1059 ( \631 , \629 , \630 );
mxor \mul_6_11/U$1055 ( \632 , \628 , \631 );
mand \mul_6_11/U$1015 ( \633 , \317_A[8] , \239_B[5] );
mxor \mul_6_11/U$970 ( \634 , \632 , \633 );
mand \mul_6_11/U$974 ( \635 , \562 , \563 );
mand \mul_6_11/U$973 ( \636 , \564 , \567 );
mor \mul_6_11/U$971 ( \637 , \635 , \636 );
mxor \mul_6_11/U$967 ( \638 , \634 , \637 );
mand \mul_6_11/U$923 ( \639 , \277_A[7] , \273_B[6] );
mxor \mul_6_11/U$882 ( \640 , \638 , \639 );
mand \mul_6_11/U$886 ( \641 , \568 , \569 );
mand \mul_6_11/U$885 ( \642 , \570 , \573 );
mor \mul_6_11/U$883 ( \643 , \641 , \642 );
mxor \mul_6_11/U$879 ( \644 , \640 , \643 );
mand \mul_6_11/U$831 ( \645 , \243_A[6] , \313_B[7] );
mxor \mul_6_11/U$794 ( \646 , \644 , \645 );
mand \mul_6_11/U$798 ( \647 , \574 , \575 );
mand \mul_6_11/U$797 ( \648 , \576 , \579 );
mor \mul_6_11/U$795 ( \649 , \647 , \648 );
mxor \mul_6_11/U$791 ( \650 , \646 , \649 );
mand \mul_6_11/U$739 ( \651 , \215_A[5] , \359_B[8] );
mxor \mul_6_11/U$706 ( \652 , \650 , \651 );
mand \mul_6_11/U$710 ( \653 , \580 , \581 );
mand \mul_6_11/U$709 ( \654 , \582 , \585 );
mor \mul_6_11/U$707 ( \655 , \653 , \654 );
mxor \mul_6_11/U$703 ( \656 , \652 , \655 );
mand \mul_6_11/U$647 ( \657 , \193_A[4] , \411_B[9] );
mxor \mul_6_11/U$618 ( \658 , \656 , \657 );
mand \mul_6_11/U$622 ( \659 , \586 , \587 );
mand \mul_6_11/U$621 ( \660 , \588 , \591 );
mor \mul_6_11/U$619 ( \661 , \659 , \660 );
mxor \mul_6_11/U$615 ( \662 , \658 , \661 );
mand \mul_6_11/U$555 ( \663 , \177_A[3] , \469_B[10] );
mxor \mul_6_11/U$530 ( \664 , \662 , \663 );
mand \mul_6_11/U$534 ( \665 , \592 , \593 );
mand \mul_6_11/U$533 ( \666 , \594 , \597 );
mor \mul_6_11/U$531 ( \667 , \665 , \666 );
mxor \mul_6_11/U$527 ( \668 , \664 , \667 );
mand \mul_6_11/U$463 ( \669 , \167_A[2] , \533_B[11] );
mxor \mul_6_11/U$442 ( \670 , \668 , \669 );
mand \mul_6_11/U$446 ( \671 , \598 , \599 );
mand \mul_6_11/U$445 ( \672 , \600 , \601 );
mor \mul_6_11/U$443 ( \673 , \671 , \672 );
mxor \mul_6_11/U$439 ( \674 , \670 , \673 );
mand \mul_6_11/U$371 ( \675 , \161_A[1] , \603_B[12] );
mxor \mul_6_11/U$354 ( \676 , \674 , \675 );
mand \mul_6_11/U$355 ( \677 , \602 , \604 );
mxor \mul_6_11/U$351 ( \678 , \676 , \677 );
mbuf \mul_6_11/B[13] ( \679_B[13] , \b[13] );
mand \mul_6_11/U$279 ( \680 , \156_A[0] , \679_B[13] );
mxor \mul_6_11/U$263 ( \681 , \678 , \680 );
mbuf \mul_6_11/Z[13] ( \682_Z[13] , \681 );
mbuf \mul_6_11/A[14] ( \683_A[14] , \a[14] );
mand \mul_6_11/U$1394 ( \684 , \683_A[14] , \157_B[0] );
mand \mul_6_11/U$1379 ( \685 , \607_A[13] , \163_B[1] );
mxor \mul_6_11/U$1314 ( \686 , \684 , \685 );
mand \mul_6_11/U$1318 ( \687 , \608 , \609 );
mand \mul_6_11/U$1317 ( \688 , \610 , \613 );
mor \mul_6_11/U$1315 ( \689 , \687 , \688 );
mxor \mul_6_11/U$1311 ( \690 , \686 , \689 );
mand \mul_6_11/U$1290 ( \691 , \537_A[12] , \173_B[2] );
mxor \mul_6_11/U$1229 ( \692 , \690 , \691 );
mand \mul_6_11/U$1233 ( \693 , \614 , \615 );
mand \mul_6_11/U$1232 ( \694 , \616 , \619 );
mor \mul_6_11/U$1230 ( \695 , \693 , \694 );
mxor \mul_6_11/U$1226 ( \696 , \692 , \695 );
mand \mul_6_11/U$1198 ( \697 , \473_A[11] , \189_B[3] );
mxor \mul_6_11/U$1141 ( \698 , \696 , \697 );
mand \mul_6_11/U$1145 ( \699 , \620 , \621 );
mand \mul_6_11/U$1144 ( \700 , \622 , \625 );
mor \mul_6_11/U$1142 ( \701 , \699 , \700 );
mxor \mul_6_11/U$1138 ( \702 , \698 , \701 );
mand \mul_6_11/U$1106 ( \703 , \415_A[10] , \211_B[4] );
mxor \mul_6_11/U$1053 ( \704 , \702 , \703 );
mand \mul_6_11/U$1057 ( \705 , \626 , \627 );
mand \mul_6_11/U$1056 ( \706 , \628 , \631 );
mor \mul_6_11/U$1054 ( \707 , \705 , \706 );
mxor \mul_6_11/U$1050 ( \708 , \704 , \707 );
mand \mul_6_11/U$1014 ( \709 , \363_A[9] , \239_B[5] );
mxor \mul_6_11/U$965 ( \710 , \708 , \709 );
mand \mul_6_11/U$969 ( \711 , \632 , \633 );
mand \mul_6_11/U$968 ( \712 , \634 , \637 );
mor \mul_6_11/U$966 ( \713 , \711 , \712 );
mxor \mul_6_11/U$962 ( \714 , \710 , \713 );
mand \mul_6_11/U$922 ( \715 , \317_A[8] , \273_B[6] );
mxor \mul_6_11/U$877 ( \716 , \714 , \715 );
mand \mul_6_11/U$881 ( \717 , \638 , \639 );
mand \mul_6_11/U$880 ( \718 , \640 , \643 );
mor \mul_6_11/U$878 ( \719 , \717 , \718 );
mxor \mul_6_11/U$874 ( \720 , \716 , \719 );
mand \mul_6_11/U$830 ( \721 , \277_A[7] , \313_B[7] );
mxor \mul_6_11/U$789 ( \722 , \720 , \721 );
mand \mul_6_11/U$793 ( \723 , \644 , \645 );
mand \mul_6_11/U$792 ( \724 , \646 , \649 );
mor \mul_6_11/U$790 ( \725 , \723 , \724 );
mxor \mul_6_11/U$786 ( \726 , \722 , \725 );
mand \mul_6_11/U$738 ( \727 , \243_A[6] , \359_B[8] );
mxor \mul_6_11/U$701 ( \728 , \726 , \727 );
mand \mul_6_11/U$705 ( \729 , \650 , \651 );
mand \mul_6_11/U$704 ( \730 , \652 , \655 );
mor \mul_6_11/U$702 ( \731 , \729 , \730 );
mxor \mul_6_11/U$698 ( \732 , \728 , \731 );
mand \mul_6_11/U$646 ( \733 , \215_A[5] , \411_B[9] );
mxor \mul_6_11/U$613 ( \734 , \732 , \733 );
mand \mul_6_11/U$617 ( \735 , \656 , \657 );
mand \mul_6_11/U$616 ( \736 , \658 , \661 );
mor \mul_6_11/U$614 ( \737 , \735 , \736 );
mxor \mul_6_11/U$610 ( \738 , \734 , \737 );
mand \mul_6_11/U$554 ( \739 , \193_A[4] , \469_B[10] );
mxor \mul_6_11/U$525 ( \740 , \738 , \739 );
mand \mul_6_11/U$529 ( \741 , \662 , \663 );
mand \mul_6_11/U$528 ( \742 , \664 , \667 );
mor \mul_6_11/U$526 ( \743 , \741 , \742 );
mxor \mul_6_11/U$522 ( \744 , \740 , \743 );
mand \mul_6_11/U$462 ( \745 , \177_A[3] , \533_B[11] );
mxor \mul_6_11/U$437 ( \746 , \744 , \745 );
mand \mul_6_11/U$441 ( \747 , \668 , \669 );
mand \mul_6_11/U$440 ( \748 , \670 , \673 );
mor \mul_6_11/U$438 ( \749 , \747 , \748 );
mxor \mul_6_11/U$434 ( \750 , \746 , \749 );
mand \mul_6_11/U$370 ( \751 , \167_A[2] , \603_B[12] );
mxor \mul_6_11/U$349 ( \752 , \750 , \751 );
mand \mul_6_11/U$353 ( \753 , \674 , \675 );
mand \mul_6_11/U$352 ( \754 , \676 , \677 );
mor \mul_6_11/U$350 ( \755 , \753 , \754 );
mxor \mul_6_11/U$346 ( \756 , \752 , \755 );
mand \mul_6_11/U$278 ( \757 , \161_A[1] , \679_B[13] );
mxor \mul_6_11/U$261 ( \758 , \756 , \757 );
mand \mul_6_11/U$262 ( \759 , \678 , \680 );
mxor \mul_6_11/U$258 ( \760 , \758 , \759 );
mbuf \mul_6_11/B[14] ( \761_B[14] , \b[14] );
mand \mul_6_11/U$186 ( \762 , \156_A[0] , \761_B[14] );
mxor \mul_6_11/U$170 ( \763 , \760 , \762 );
mbuf \mul_6_11/Z[14] ( \764_Z[14] , \763 );
mbuf \mul_6_11/A[15] ( \765_A[15] , \a[15] );
mand \mul_6_11/U$1393 ( \766 , \765_A[15] , \157_B[0] );
mand \mul_6_11/U$1378 ( \767 , \683_A[14] , \163_B[1] );
mxor \mul_6_11/U$1309 ( \768 , \766 , \767 );
mand \mul_6_11/U$1313 ( \769 , \684 , \685 );
mand \mul_6_11/U$1312 ( \770 , \686 , \689 );
mor \mul_6_11/U$1310 ( \771 , \769 , \770 );
mxor \mul_6_11/U$1306 ( \772 , \768 , \771 );
mand \mul_6_11/U$1289 ( \773 , \607_A[13] , \173_B[2] );
mxor \mul_6_11/U$1224 ( \774 , \772 , \773 );
mand \mul_6_11/U$1228 ( \775 , \690 , \691 );
mand \mul_6_11/U$1227 ( \776 , \692 , \695 );
mor \mul_6_11/U$1225 ( \777 , \775 , \776 );
mxor \mul_6_11/U$1221 ( \778 , \774 , \777 );
mand \mul_6_11/U$1197 ( \779 , \537_A[12] , \189_B[3] );
mxor \mul_6_11/U$1136 ( \780 , \778 , \779 );
mand \mul_6_11/U$1140 ( \781 , \696 , \697 );
mand \mul_6_11/U$1139 ( \782 , \698 , \701 );
mor \mul_6_11/U$1137 ( \783 , \781 , \782 );
mxor \mul_6_11/U$1133 ( \784 , \780 , \783 );
mand \mul_6_11/U$1105 ( \785 , \473_A[11] , \211_B[4] );
mxor \mul_6_11/U$1048 ( \786 , \784 , \785 );
mand \mul_6_11/U$1052 ( \787 , \702 , \703 );
mand \mul_6_11/U$1051 ( \788 , \704 , \707 );
mor \mul_6_11/U$1049 ( \789 , \787 , \788 );
mxor \mul_6_11/U$1045 ( \790 , \786 , \789 );
mand \mul_6_11/U$1013 ( \791 , \415_A[10] , \239_B[5] );
mxor \mul_6_11/U$960 ( \792 , \790 , \791 );
mand \mul_6_11/U$964 ( \793 , \708 , \709 );
mand \mul_6_11/U$963 ( \794 , \710 , \713 );
mor \mul_6_11/U$961 ( \795 , \793 , \794 );
mxor \mul_6_11/U$957 ( \796 , \792 , \795 );
mand \mul_6_11/U$921 ( \797 , \363_A[9] , \273_B[6] );
mxor \mul_6_11/U$872 ( \798 , \796 , \797 );
mand \mul_6_11/U$876 ( \799 , \714 , \715 );
mand \mul_6_11/U$875 ( \800 , \716 , \719 );
mor \mul_6_11/U$873 ( \801 , \799 , \800 );
mxor \mul_6_11/U$869 ( \802 , \798 , \801 );
mand \mul_6_11/U$829 ( \803 , \317_A[8] , \313_B[7] );
mxor \mul_6_11/U$784 ( \804 , \802 , \803 );
mand \mul_6_11/U$788 ( \805 , \720 , \721 );
mand \mul_6_11/U$787 ( \806 , \722 , \725 );
mor \mul_6_11/U$785 ( \807 , \805 , \806 );
mxor \mul_6_11/U$781 ( \808 , \804 , \807 );
mand \mul_6_11/U$737 ( \809 , \277_A[7] , \359_B[8] );
mxor \mul_6_11/U$696 ( \810 , \808 , \809 );
mand \mul_6_11/U$700 ( \811 , \726 , \727 );
mand \mul_6_11/U$699 ( \812 , \728 , \731 );
mor \mul_6_11/U$697 ( \813 , \811 , \812 );
mxor \mul_6_11/U$693 ( \814 , \810 , \813 );
mand \mul_6_11/U$645 ( \815 , \243_A[6] , \411_B[9] );
mxor \mul_6_11/U$608 ( \816 , \814 , \815 );
mand \mul_6_11/U$612 ( \817 , \732 , \733 );
mand \mul_6_11/U$611 ( \818 , \734 , \737 );
mor \mul_6_11/U$609 ( \819 , \817 , \818 );
mxor \mul_6_11/U$605 ( \820 , \816 , \819 );
mand \mul_6_11/U$553 ( \821 , \215_A[5] , \469_B[10] );
mxor \mul_6_11/U$520 ( \822 , \820 , \821 );
mand \mul_6_11/U$524 ( \823 , \738 , \739 );
mand \mul_6_11/U$523 ( \824 , \740 , \743 );
mor \mul_6_11/U$521 ( \825 , \823 , \824 );
mxor \mul_6_11/U$517 ( \826 , \822 , \825 );
mand \mul_6_11/U$461 ( \827 , \193_A[4] , \533_B[11] );
mxor \mul_6_11/U$432 ( \828 , \826 , \827 );
mand \mul_6_11/U$436 ( \829 , \744 , \745 );
mand \mul_6_11/U$435 ( \830 , \746 , \749 );
mor \mul_6_11/U$433 ( \831 , \829 , \830 );
mxor \mul_6_11/U$429 ( \832 , \828 , \831 );
mand \mul_6_11/U$369 ( \833 , \177_A[3] , \603_B[12] );
mxor \mul_6_11/U$344 ( \834 , \832 , \833 );
mand \mul_6_11/U$348 ( \835 , \750 , \751 );
mand \mul_6_11/U$347 ( \836 , \752 , \755 );
mor \mul_6_11/U$345 ( \837 , \835 , \836 );
mxor \mul_6_11/U$341 ( \838 , \834 , \837 );
mand \mul_6_11/U$277 ( \839 , \167_A[2] , \679_B[13] );
mxor \mul_6_11/U$256 ( \840 , \838 , \839 );
mand \mul_6_11/U$260 ( \841 , \756 , \757 );
mand \mul_6_11/U$259 ( \842 , \758 , \759 );
mor \mul_6_11/U$257 ( \843 , \841 , \842 );
mxor \mul_6_11/U$253 ( \844 , \840 , \843 );
mand \mul_6_11/U$185 ( \845 , \161_A[1] , \761_B[14] );
mxor \mul_6_11/U$168 ( \846 , \844 , \845 );
mand \mul_6_11/U$169 ( \847 , \760 , \762 );
mxor \mul_6_11/U$165 ( \848 , \846 , \847 );
mbuf \mul_6_11/B[15] ( \849_B[15] , \b[15] );
mand \mul_6_11/U$93 ( \850 , \156_A[0] , \849_B[15] );
mxor \mul_6_11/U$77 ( \851 , \848 , \850 );
mbuf \mul_6_11/Z[15] ( \852_Z[15] , \851 );
mnor \U$10 ( \853 , \160 , \166_Z[1] , \176_Z[2] , \192_Z[3] , \214_Z[4] , \242_Z[5] , \276_Z[6] , \316_Z[7] , \362_Z[8] , \414_Z[9] , \472_Z[10] , \536_Z[11] , \606_Z[12] , \682_Z[13] , \764_Z[14] , \852_Z[15] );
mnot \U$7 ( \854 , \166_Z[1] );
mnor \U$8 ( \855 , \159_Z[0] , \854 , \176_Z[2] , \192_Z[3] , \214_Z[4] , \242_Z[5] , \276_Z[6] , \316_Z[7] , \362_Z[8] , \414_Z[9] , \472_Z[10] , \536_Z[11] , \606_Z[12] , \682_Z[13] , \764_Z[14] , \852_Z[15] );
mnot \U$11 ( \856 , \176_Z[2] );
mnor \U$12 ( \857 , \159_Z[0] , \166_Z[1] , \856 , \192_Z[3] , \214_Z[4] , \242_Z[5] , \276_Z[6] , \316_Z[7] , \362_Z[8] , \414_Z[9] , \472_Z[10] , \536_Z[11] , \606_Z[12] , \682_Z[13] , \764_Z[14] , \852_Z[15] );
mnot \U$13 ( \858 , \192_Z[3] );
mnor \U$14 ( \859 , \159_Z[0] , \166_Z[1] , \176_Z[2] , \858 , \214_Z[4] , \242_Z[5] , \276_Z[6] , \316_Z[7] , \362_Z[8] , \414_Z[9] , \472_Z[10] , \536_Z[11] , \606_Z[12] , \682_Z[13] , \764_Z[14] , \852_Z[15] );
mnot \U$15 ( \860 , \214_Z[4] );
mnor \U$16 ( \861 , \159_Z[0] , \166_Z[1] , \176_Z[2] , \192_Z[3] , \860 , \242_Z[5] , \276_Z[6] , \316_Z[7] , \362_Z[8] , \414_Z[9] , \472_Z[10] , \536_Z[11] , \606_Z[12] , \682_Z[13] , \764_Z[14] , \852_Z[15] );
mnot \U$17 ( \862 , \242_Z[5] );
mnor \U$18 ( \863 , \159_Z[0] , \166_Z[1] , \176_Z[2] , \192_Z[3] , \214_Z[4] , \862 , \276_Z[6] , \316_Z[7] , \362_Z[8] , \414_Z[9] , \472_Z[10] , \536_Z[11] , \606_Z[12] , \682_Z[13] , \764_Z[14] , \852_Z[15] );
mnot \U$19 ( \864 , \276_Z[6] );
mnor \U$20 ( \865 , \159_Z[0] , \166_Z[1] , \176_Z[2] , \192_Z[3] , \214_Z[4] , \242_Z[5] , \864 , \316_Z[7] , \362_Z[8] , \414_Z[9] , \472_Z[10] , \536_Z[11] , \606_Z[12] , \682_Z[13] , \764_Z[14] , \852_Z[15] );
mnot \U$21 ( \866 , \316_Z[7] );
mnor \U$22 ( \867 , \159_Z[0] , \166_Z[1] , \176_Z[2] , \192_Z[3] , \214_Z[4] , \242_Z[5] , \276_Z[6] , \866 , \362_Z[8] , \414_Z[9] , \472_Z[10] , \536_Z[11] , \606_Z[12] , \682_Z[13] , \764_Z[14] , \852_Z[15] );
mnot \U$23 ( \868 , \362_Z[8] );
mnor \U$24 ( \869 , \159_Z[0] , \166_Z[1] , \176_Z[2] , \192_Z[3] , \214_Z[4] , \242_Z[5] , \276_Z[6] , \316_Z[7] , \868 , \414_Z[9] , \472_Z[10] , \536_Z[11] , \606_Z[12] , \682_Z[13] , \764_Z[14] , \852_Z[15] );
mnot \U$25 ( \870 , \414_Z[9] );
mnor \U$26 ( \871 , \159_Z[0] , \166_Z[1] , \176_Z[2] , \192_Z[3] , \214_Z[4] , \242_Z[5] , \276_Z[6] , \316_Z[7] , \362_Z[8] , \870 , \472_Z[10] , \536_Z[11] , \606_Z[12] , \682_Z[13] , \764_Z[14] , \852_Z[15] );
mnot \U$27 ( \872 , \472_Z[10] );
mnor \U$28 ( \873 , \159_Z[0] , \166_Z[1] , \176_Z[2] , \192_Z[3] , \214_Z[4] , \242_Z[5] , \276_Z[6] , \316_Z[7] , \362_Z[8] , \414_Z[9] , \872 , \536_Z[11] , \606_Z[12] , \682_Z[13] , \764_Z[14] , \852_Z[15] );
mnot \U$29 ( \874 , \536_Z[11] );
mnor \U$30 ( \875 , \159_Z[0] , \166_Z[1] , \176_Z[2] , \192_Z[3] , \214_Z[4] , \242_Z[5] , \276_Z[6] , \316_Z[7] , \362_Z[8] , \414_Z[9] , \472_Z[10] , \874 , \606_Z[12] , \682_Z[13] , \764_Z[14] , \852_Z[15] );
mnor \U$6 ( \876 , \853 , \855 , \857 , \859 , \861 , \863 , \865 , \867 , \869 , \871 , \873 , \875 );
m_DC \n22[0]_g1 ( \877 , 1'b0 , \876 );
mor \U$5/U$1 ( \878 , \a[0] , \d[0] );
mand \U$1/U$13 ( \879 , \878 , \875 );
mand \U$4/U$1 ( \880 , \b[0] , \c[0] );
mand \U$1/U$12 ( \881 , \880 , \873 );
mor \U$3/U$1 ( \882 , \a[0] , \b[0] );
mand \U$1/U$11 ( \883 , \882 , \871 );
mxor \U$2/U$1 ( \884 , \c[0] , \d[0] );
mand \U$1/U$10 ( \885 , \884 , \869 );
mbuf \mul_17_13/A[0] ( \886_A[0] , \b[0] );
mbuf \mul_17_13/B[0] ( \887_B[0] , \c[0] );
mand \mul_17_13/U$1408 ( \888 , \886_A[0] , \887_B[0] );
mbuf \mul_17_13/Z[0] ( \889_Z[0] , \888 );
mand \U$1/U$9 ( \890 , \889_Z[0] , \867 );
mbuf \mul_16_12/A[0] ( \891_A[0] , \a[0] );
mbuf \mul_16_12/B[0] ( \892_B[0] , \d[0] );
mand \mul_16_12/U$1408 ( \893 , \891_A[0] , \892_B[0] );
mbuf \mul_16_12/Z[0] ( \894_Z[0] , \893 );
mand \U$1/U$8 ( \895 , \894_Z[0] , \865 );
mbuf \add_15_12/A[0] ( \896_A[0] , \b[0] );
mbuf \add_15_12/B[0] ( \897_B[0] , \d[0] );
mxor \add_15_12/U$88 ( \898 , \896_A[0] , \897_B[0] );
mbuf \add_15_12/SUM[0] ( \899_SUM[0] , \898 );
mand \U$1/U$7 ( \900 , \899_SUM[0] , \863 );
mbuf \add_14_12/A[0] ( \901_A[0] , \a[0] );
mbuf \add_14_12/B[0] ( \902_B[0] , \c[0] );
mxor \add_14_12/U$88 ( \903 , \901_A[0] , \902_B[0] );
mbuf \add_14_12/SUM[0] ( \904_SUM[0] , \903 );
mand \U$1/U$6 ( \905 , \904_SUM[0] , \861 );
mand \U$1/U$5 ( \906 , \d[0] , \859 );
mand \U$1/U$4 ( \907 , \c[0] , \857 );
mand \U$1/U$3 ( \908 , \b[0] , \855 );
mand \U$1/U$2 ( \909 , \a[0] , \853 );
mor \U$1/U$1 ( \910 , \877 , \879 , \881 , \883 , \885 , \890 , \895 , \900 , \905 , \906 , \907 , \908 , \909 );
m_DC \n22[1]_g1 ( \911 , 1'b0 , \876 );
mor \U$5/U$2 ( \912 , \a[1] , \d[1] );
mand \U$1/U$27 ( \913 , \912 , \875 );
mand \U$4/U$2 ( \914 , \b[1] , \c[1] );
mand \U$1/U$26 ( \915 , \914 , \873 );
mor \U$3/U$2 ( \916 , \a[1] , \b[1] );
mand \U$1/U$25 ( \917 , \916 , \871 );
mxor \U$2/U$2 ( \918 , \c[1] , \d[1] );
mand \U$1/U$24 ( \919 , \918 , \869 );
mbuf \mul_17_13/A[1] ( \920_A[1] , \b[1] );
mand \mul_17_13/U$1407 ( \921 , \920_A[1] , \887_B[0] );
mbuf \mul_17_13/B[1] ( \922_B[1] , \c[1] );
mand \mul_17_13/U$1392 ( \923 , \886_A[0] , \922_B[1] );
mxor \mul_17_13/U$1376 ( \924 , \921 , \923 );
mbuf \mul_17_13/Z[1] ( \925_Z[1] , \924 );
mand \U$1/U$23 ( \926 , \925_Z[1] , \867 );
mbuf \mul_16_12/A[1] ( \927_A[1] , \a[1] );
mand \mul_16_12/U$1407 ( \928 , \927_A[1] , \892_B[0] );
mbuf \mul_16_12/B[1] ( \929_B[1] , \d[1] );
mand \mul_16_12/U$1392 ( \930 , \891_A[0] , \929_B[1] );
mxor \mul_16_12/U$1376 ( \931 , \928 , \930 );
mbuf \mul_16_12/Z[1] ( \932_Z[1] , \931 );
mand \U$1/U$22 ( \933 , \932_Z[1] , \865 );
mbuf \add_15_12/A[1] ( \934_A[1] , \b[1] );
mbuf \add_15_12/B[1] ( \935_B[1] , \d[1] );
mxor \add_15_12/U$86 ( \936 , \934_A[1] , \935_B[1] );
mand \add_15_12/U$87 ( \937 , \896_A[0] , \897_B[0] );
mxor \add_15_12/U$85 ( \938 , \936 , \937 );
mbuf \add_15_12/SUM[1] ( \939_SUM[1] , \938 );
mand \U$1/U$21 ( \940 , \939_SUM[1] , \863 );
mbuf \add_14_12/A[1] ( \941_A[1] , \a[1] );
mbuf \add_14_12/B[1] ( \942_B[1] , \c[1] );
mxor \add_14_12/U$86 ( \943 , \941_A[1] , \942_B[1] );
mand \add_14_12/U$87 ( \944 , \901_A[0] , \902_B[0] );
mxor \add_14_12/U$85 ( \945 , \943 , \944 );
mbuf \add_14_12/SUM[1] ( \946_SUM[1] , \945 );
mand \U$1/U$20 ( \947 , \946_SUM[1] , \861 );
mand \U$1/U$19 ( \948 , \d[1] , \859 );
mand \U$1/U$18 ( \949 , \c[1] , \857 );
mand \U$1/U$17 ( \950 , \b[1] , \855 );
mand \U$1/U$16 ( \951 , \a[1] , \853 );
mor \U$1/U$15 ( \952 , \911 , \913 , \915 , \917 , \919 , \926 , \933 , \940 , \947 , \948 , \949 , \950 , \951 );
m_DC \n22[2]_g1 ( \953 , 1'b0 , \876 );
mor \U$5/U$3 ( \954 , \a[2] , \d[2] );
mand \U$1/U$41 ( \955 , \954 , \875 );
mand \U$4/U$3 ( \956 , \b[2] , \c[2] );
mand \U$1/U$40 ( \957 , \956 , \873 );
mor \U$3/U$3 ( \958 , \a[2] , \b[2] );
mand \U$1/U$39 ( \959 , \958 , \871 );
mxor \U$2/U$3 ( \960 , \c[2] , \d[2] );
mand \U$1/U$38 ( \961 , \960 , \869 );
mbuf \mul_17_13/A[2] ( \962_A[2] , \b[2] );
mand \mul_17_13/U$1406 ( \963 , \962_A[2] , \887_B[0] );
mand \mul_17_13/U$1391 ( \964 , \920_A[1] , \922_B[1] );
mxor \mul_17_13/U$1374 ( \965 , \963 , \964 );
mand \mul_17_13/U$1375 ( \966 , \921 , \923 );
mxor \mul_17_13/U$1371 ( \967 , \965 , \966 );
mbuf \mul_17_13/B[2] ( \968_B[2] , \c[2] );
mand \mul_17_13/U$1302 ( \969 , \886_A[0] , \968_B[2] );
mxor \mul_17_13/U$1286 ( \970 , \967 , \969 );
mbuf \mul_17_13/Z[2] ( \971_Z[2] , \970 );
mand \U$1/U$37 ( \972 , \971_Z[2] , \867 );
mbuf \mul_16_12/A[2] ( \973_A[2] , \a[2] );
mand \mul_16_12/U$1406 ( \974 , \973_A[2] , \892_B[0] );
mand \mul_16_12/U$1391 ( \975 , \927_A[1] , \929_B[1] );
mxor \mul_16_12/U$1374 ( \976 , \974 , \975 );
mand \mul_16_12/U$1375 ( \977 , \928 , \930 );
mxor \mul_16_12/U$1371 ( \978 , \976 , \977 );
mbuf \mul_16_12/B[2] ( \979_B[2] , \d[2] );
mand \mul_16_12/U$1302 ( \980 , \891_A[0] , \979_B[2] );
mxor \mul_16_12/U$1286 ( \981 , \978 , \980 );
mbuf \mul_16_12/Z[2] ( \982_Z[2] , \981 );
mand \U$1/U$36 ( \983 , \982_Z[2] , \865 );
mbuf \add_15_12/A[2] ( \984_A[2] , \b[2] );
mbuf \add_15_12/B[2] ( \985_B[2] , \d[2] );
mxor \add_15_12/U$80 ( \986 , \984_A[2] , \985_B[2] );
mand \add_15_12/U$84 ( \987 , \934_A[1] , \935_B[1] );
mand \add_15_12/U$83 ( \988 , \935_B[1] , \937 );
mand \add_15_12/U$82 ( \989 , \934_A[1] , \937 );
mor \add_15_12/U$81 ( \990 , \987 , \988 , \989 );
mxor \add_15_12/U$79 ( \991 , \986 , \990 );
mbuf \add_15_12/SUM[2] ( \992_SUM[2] , \991 );
mand \U$1/U$35 ( \993 , \992_SUM[2] , \863 );
mbuf \add_14_12/A[2] ( \994_A[2] , \a[2] );
mbuf \add_14_12/B[2] ( \995_B[2] , \c[2] );
mxor \add_14_12/U$80 ( \996 , \994_A[2] , \995_B[2] );
mand \add_14_12/U$84 ( \997 , \941_A[1] , \942_B[1] );
mand \add_14_12/U$83 ( \998 , \942_B[1] , \944 );
mand \add_14_12/U$82 ( \999 , \941_A[1] , \944 );
mor \add_14_12/U$81 ( \1000 , \997 , \998 , \999 );
mxor \add_14_12/U$79 ( \1001 , \996 , \1000 );
mbuf \add_14_12/SUM[2] ( \1002_SUM[2] , \1001 );
mand \U$1/U$34 ( \1003 , \1002_SUM[2] , \861 );
mand \U$1/U$33 ( \1004 , \d[2] , \859 );
mand \U$1/U$32 ( \1005 , \c[2] , \857 );
mand \U$1/U$31 ( \1006 , \b[2] , \855 );
mand \U$1/U$30 ( \1007 , \a[2] , \853 );
mor \U$1/U$29 ( \1008 , \953 , \955 , \957 , \959 , \961 , \972 , \983 , \993 , \1003 , \1004 , \1005 , \1006 , \1007 );
m_DC \n22[3]_g1 ( \1009 , 1'b0 , \876 );
mor \U$5/U$4 ( \1010 , \a[3] , \d[3] );
mand \U$1/U$55 ( \1011 , \1010 , \875 );
mand \U$4/U$4 ( \1012 , \b[3] , \c[3] );
mand \U$1/U$54 ( \1013 , \1012 , \873 );
mor \U$3/U$4 ( \1014 , \a[3] , \b[3] );
mand \U$1/U$53 ( \1015 , \1014 , \871 );
mxor \U$2/U$4 ( \1016 , \c[3] , \d[3] );
mand \U$1/U$52 ( \1017 , \1016 , \869 );
mbuf \mul_17_13/A[3] ( \1018_A[3] , \b[3] );
mand \mul_17_13/U$1405 ( \1019 , \1018_A[3] , \887_B[0] );
mand \mul_17_13/U$1390 ( \1020 , \962_A[2] , \922_B[1] );
mxor \mul_17_13/U$1369 ( \1021 , \1019 , \1020 );
mand \mul_17_13/U$1373 ( \1022 , \963 , \964 );
mand \mul_17_13/U$1372 ( \1023 , \965 , \966 );
mor \mul_17_13/U$1370 ( \1024 , \1022 , \1023 );
mxor \mul_17_13/U$1366 ( \1025 , \1021 , \1024 );
mand \mul_17_13/U$1301 ( \1026 , \920_A[1] , \968_B[2] );
mxor \mul_17_13/U$1284 ( \1027 , \1025 , \1026 );
mand \mul_17_13/U$1285 ( \1028 , \967 , \969 );
mxor \mul_17_13/U$1281 ( \1029 , \1027 , \1028 );
mbuf \mul_17_13/B[3] ( \1030_B[3] , \c[3] );
mand \mul_17_13/U$1209 ( \1031 , \886_A[0] , \1030_B[3] );
mxor \mul_17_13/U$1193 ( \1032 , \1029 , \1031 );
mbuf \mul_17_13/Z[3] ( \1033_Z[3] , \1032 );
mand \U$1/U$51 ( \1034 , \1033_Z[3] , \867 );
mbuf \mul_16_12/A[3] ( \1035_A[3] , \a[3] );
mand \mul_16_12/U$1405 ( \1036 , \1035_A[3] , \892_B[0] );
mand \mul_16_12/U$1390 ( \1037 , \973_A[2] , \929_B[1] );
mxor \mul_16_12/U$1369 ( \1038 , \1036 , \1037 );
mand \mul_16_12/U$1373 ( \1039 , \974 , \975 );
mand \mul_16_12/U$1372 ( \1040 , \976 , \977 );
mor \mul_16_12/U$1370 ( \1041 , \1039 , \1040 );
mxor \mul_16_12/U$1366 ( \1042 , \1038 , \1041 );
mand \mul_16_12/U$1301 ( \1043 , \927_A[1] , \979_B[2] );
mxor \mul_16_12/U$1284 ( \1044 , \1042 , \1043 );
mand \mul_16_12/U$1285 ( \1045 , \978 , \980 );
mxor \mul_16_12/U$1281 ( \1046 , \1044 , \1045 );
mbuf \mul_16_12/B[3] ( \1047_B[3] , \d[3] );
mand \mul_16_12/U$1209 ( \1048 , \891_A[0] , \1047_B[3] );
mxor \mul_16_12/U$1193 ( \1049 , \1046 , \1048 );
mbuf \mul_16_12/Z[3] ( \1050_Z[3] , \1049 );
mand \U$1/U$50 ( \1051 , \1050_Z[3] , \865 );
mbuf \add_15_12/A[3] ( \1052_A[3] , \b[3] );
mbuf \add_15_12/B[3] ( \1053_B[3] , \d[3] );
mxor \add_15_12/U$74 ( \1054 , \1052_A[3] , \1053_B[3] );
mand \add_15_12/U$78 ( \1055 , \984_A[2] , \985_B[2] );
mand \add_15_12/U$77 ( \1056 , \985_B[2] , \990 );
mand \add_15_12/U$76 ( \1057 , \984_A[2] , \990 );
mor \add_15_12/U$75 ( \1058 , \1055 , \1056 , \1057 );
mxor \add_15_12/U$73 ( \1059 , \1054 , \1058 );
mbuf \add_15_12/SUM[3] ( \1060_SUM[3] , \1059 );
mand \U$1/U$49 ( \1061 , \1060_SUM[3] , \863 );
mbuf \add_14_12/A[3] ( \1062_A[3] , \a[3] );
mbuf \add_14_12/B[3] ( \1063_B[3] , \c[3] );
mxor \add_14_12/U$74 ( \1064 , \1062_A[3] , \1063_B[3] );
mand \add_14_12/U$78 ( \1065 , \994_A[2] , \995_B[2] );
mand \add_14_12/U$77 ( \1066 , \995_B[2] , \1000 );
mand \add_14_12/U$76 ( \1067 , \994_A[2] , \1000 );
mor \add_14_12/U$75 ( \1068 , \1065 , \1066 , \1067 );
mxor \add_14_12/U$73 ( \1069 , \1064 , \1068 );
mbuf \add_14_12/SUM[3] ( \1070_SUM[3] , \1069 );
mand \U$1/U$48 ( \1071 , \1070_SUM[3] , \861 );
mand \U$1/U$47 ( \1072 , \d[3] , \859 );
mand \U$1/U$46 ( \1073 , \c[3] , \857 );
mand \U$1/U$45 ( \1074 , \b[3] , \855 );
mand \U$1/U$44 ( \1075 , \a[3] , \853 );
mor \U$1/U$43 ( \1076 , \1009 , \1011 , \1013 , \1015 , \1017 , \1034 , \1051 , \1061 , \1071 , \1072 , \1073 , \1074 , \1075 );
m_DC \n22[4]_g1 ( \1077 , 1'b0 , \876 );
mor \U$5/U$5 ( \1078 , \a[4] , \d[4] );
mand \U$1/U$69 ( \1079 , \1078 , \875 );
mand \U$4/U$5 ( \1080 , \b[4] , \c[4] );
mand \U$1/U$68 ( \1081 , \1080 , \873 );
mor \U$3/U$5 ( \1082 , \a[4] , \b[4] );
mand \U$1/U$67 ( \1083 , \1082 , \871 );
mxor \U$2/U$5 ( \1084 , \c[4] , \d[4] );
mand \U$1/U$66 ( \1085 , \1084 , \869 );
mbuf \mul_17_13/A[4] ( \1086_A[4] , \b[4] );
mand \mul_17_13/U$1404 ( \1087 , \1086_A[4] , \887_B[0] );
mand \mul_17_13/U$1389 ( \1088 , \1018_A[3] , \922_B[1] );
mxor \mul_17_13/U$1364 ( \1089 , \1087 , \1088 );
mand \mul_17_13/U$1368 ( \1090 , \1019 , \1020 );
mand \mul_17_13/U$1367 ( \1091 , \1021 , \1024 );
mor \mul_17_13/U$1365 ( \1092 , \1090 , \1091 );
mxor \mul_17_13/U$1361 ( \1093 , \1089 , \1092 );
mand \mul_17_13/U$1300 ( \1094 , \962_A[2] , \968_B[2] );
mxor \mul_17_13/U$1279 ( \1095 , \1093 , \1094 );
mand \mul_17_13/U$1283 ( \1096 , \1025 , \1026 );
mand \mul_17_13/U$1282 ( \1097 , \1027 , \1028 );
mor \mul_17_13/U$1280 ( \1098 , \1096 , \1097 );
mxor \mul_17_13/U$1276 ( \1099 , \1095 , \1098 );
mand \mul_17_13/U$1208 ( \1100 , \920_A[1] , \1030_B[3] );
mxor \mul_17_13/U$1191 ( \1101 , \1099 , \1100 );
mand \mul_17_13/U$1192 ( \1102 , \1029 , \1031 );
mxor \mul_17_13/U$1188 ( \1103 , \1101 , \1102 );
mbuf \mul_17_13/B[4] ( \1104_B[4] , \c[4] );
mand \mul_17_13/U$1116 ( \1105 , \886_A[0] , \1104_B[4] );
mxor \mul_17_13/U$1100 ( \1106 , \1103 , \1105 );
mbuf \mul_17_13/Z[4] ( \1107_Z[4] , \1106 );
mand \U$1/U$65 ( \1108 , \1107_Z[4] , \867 );
mbuf \mul_16_12/A[4] ( \1109_A[4] , \a[4] );
mand \mul_16_12/U$1404 ( \1110 , \1109_A[4] , \892_B[0] );
mand \mul_16_12/U$1389 ( \1111 , \1035_A[3] , \929_B[1] );
mxor \mul_16_12/U$1364 ( \1112 , \1110 , \1111 );
mand \mul_16_12/U$1368 ( \1113 , \1036 , \1037 );
mand \mul_16_12/U$1367 ( \1114 , \1038 , \1041 );
mor \mul_16_12/U$1365 ( \1115 , \1113 , \1114 );
mxor \mul_16_12/U$1361 ( \1116 , \1112 , \1115 );
mand \mul_16_12/U$1300 ( \1117 , \973_A[2] , \979_B[2] );
mxor \mul_16_12/U$1279 ( \1118 , \1116 , \1117 );
mand \mul_16_12/U$1283 ( \1119 , \1042 , \1043 );
mand \mul_16_12/U$1282 ( \1120 , \1044 , \1045 );
mor \mul_16_12/U$1280 ( \1121 , \1119 , \1120 );
mxor \mul_16_12/U$1276 ( \1122 , \1118 , \1121 );
mand \mul_16_12/U$1208 ( \1123 , \927_A[1] , \1047_B[3] );
mxor \mul_16_12/U$1191 ( \1124 , \1122 , \1123 );
mand \mul_16_12/U$1192 ( \1125 , \1046 , \1048 );
mxor \mul_16_12/U$1188 ( \1126 , \1124 , \1125 );
mbuf \mul_16_12/B[4] ( \1127_B[4] , \d[4] );
mand \mul_16_12/U$1116 ( \1128 , \891_A[0] , \1127_B[4] );
mxor \mul_16_12/U$1100 ( \1129 , \1126 , \1128 );
mbuf \mul_16_12/Z[4] ( \1130_Z[4] , \1129 );
mand \U$1/U$64 ( \1131 , \1130_Z[4] , \865 );
mbuf \add_15_12/A[4] ( \1132_A[4] , \b[4] );
mbuf \add_15_12/B[4] ( \1133_B[4] , \d[4] );
mxor \add_15_12/U$68 ( \1134 , \1132_A[4] , \1133_B[4] );
mand \add_15_12/U$72 ( \1135 , \1052_A[3] , \1053_B[3] );
mand \add_15_12/U$71 ( \1136 , \1053_B[3] , \1058 );
mand \add_15_12/U$70 ( \1137 , \1052_A[3] , \1058 );
mor \add_15_12/U$69 ( \1138 , \1135 , \1136 , \1137 );
mxor \add_15_12/U$67 ( \1139 , \1134 , \1138 );
mbuf \add_15_12/SUM[4] ( \1140_SUM[4] , \1139 );
mand \U$1/U$63 ( \1141 , \1140_SUM[4] , \863 );
mbuf \add_14_12/A[4] ( \1142_A[4] , \a[4] );
mbuf \add_14_12/B[4] ( \1143_B[4] , \c[4] );
mxor \add_14_12/U$68 ( \1144 , \1142_A[4] , \1143_B[4] );
mand \add_14_12/U$72 ( \1145 , \1062_A[3] , \1063_B[3] );
mand \add_14_12/U$71 ( \1146 , \1063_B[3] , \1068 );
mand \add_14_12/U$70 ( \1147 , \1062_A[3] , \1068 );
mor \add_14_12/U$69 ( \1148 , \1145 , \1146 , \1147 );
mxor \add_14_12/U$67 ( \1149 , \1144 , \1148 );
mbuf \add_14_12/SUM[4] ( \1150_SUM[4] , \1149 );
mand \U$1/U$62 ( \1151 , \1150_SUM[4] , \861 );
mand \U$1/U$61 ( \1152 , \d[4] , \859 );
mand \U$1/U$60 ( \1153 , \c[4] , \857 );
mand \U$1/U$59 ( \1154 , \b[4] , \855 );
mand \U$1/U$58 ( \1155 , \a[4] , \853 );
mor \U$1/U$57 ( \1156 , \1077 , \1079 , \1081 , \1083 , \1085 , \1108 , \1131 , \1141 , \1151 , \1152 , \1153 , \1154 , \1155 );
m_DC \n22[5]_g1 ( \1157 , 1'b0 , \876 );
mor \U$5/U$6 ( \1158 , \a[5] , \d[5] );
mand \U$1/U$83 ( \1159 , \1158 , \875 );
mand \U$4/U$6 ( \1160 , \b[5] , \c[5] );
mand \U$1/U$82 ( \1161 , \1160 , \873 );
mor \U$3/U$6 ( \1162 , \a[5] , \b[5] );
mand \U$1/U$81 ( \1163 , \1162 , \871 );
mxor \U$2/U$6 ( \1164 , \c[5] , \d[5] );
mand \U$1/U$80 ( \1165 , \1164 , \869 );
mbuf \mul_17_13/A[5] ( \1166_A[5] , \b[5] );
mand \mul_17_13/U$1403 ( \1167 , \1166_A[5] , \887_B[0] );
mand \mul_17_13/U$1388 ( \1168 , \1086_A[4] , \922_B[1] );
mxor \mul_17_13/U$1359 ( \1169 , \1167 , \1168 );
mand \mul_17_13/U$1363 ( \1170 , \1087 , \1088 );
mand \mul_17_13/U$1362 ( \1171 , \1089 , \1092 );
mor \mul_17_13/U$1360 ( \1172 , \1170 , \1171 );
mxor \mul_17_13/U$1356 ( \1173 , \1169 , \1172 );
mand \mul_17_13/U$1299 ( \1174 , \1018_A[3] , \968_B[2] );
mxor \mul_17_13/U$1274 ( \1175 , \1173 , \1174 );
mand \mul_17_13/U$1278 ( \1176 , \1093 , \1094 );
mand \mul_17_13/U$1277 ( \1177 , \1095 , \1098 );
mor \mul_17_13/U$1275 ( \1178 , \1176 , \1177 );
mxor \mul_17_13/U$1271 ( \1179 , \1175 , \1178 );
mand \mul_17_13/U$1207 ( \1180 , \962_A[2] , \1030_B[3] );
mxor \mul_17_13/U$1186 ( \1181 , \1179 , \1180 );
mand \mul_17_13/U$1190 ( \1182 , \1099 , \1100 );
mand \mul_17_13/U$1189 ( \1183 , \1101 , \1102 );
mor \mul_17_13/U$1187 ( \1184 , \1182 , \1183 );
mxor \mul_17_13/U$1183 ( \1185 , \1181 , \1184 );
mand \mul_17_13/U$1115 ( \1186 , \920_A[1] , \1104_B[4] );
mxor \mul_17_13/U$1098 ( \1187 , \1185 , \1186 );
mand \mul_17_13/U$1099 ( \1188 , \1103 , \1105 );
mxor \mul_17_13/U$1095 ( \1189 , \1187 , \1188 );
mbuf \mul_17_13/B[5] ( \1190_B[5] , \c[5] );
mand \mul_17_13/U$1023 ( \1191 , \886_A[0] , \1190_B[5] );
mxor \mul_17_13/U$1007 ( \1192 , \1189 , \1191 );
mbuf \mul_17_13/Z[5] ( \1193_Z[5] , \1192 );
mand \U$1/U$79 ( \1194 , \1193_Z[5] , \867 );
mbuf \mul_16_12/A[5] ( \1195_A[5] , \a[5] );
mand \mul_16_12/U$1403 ( \1196 , \1195_A[5] , \892_B[0] );
mand \mul_16_12/U$1388 ( \1197 , \1109_A[4] , \929_B[1] );
mxor \mul_16_12/U$1359 ( \1198 , \1196 , \1197 );
mand \mul_16_12/U$1363 ( \1199 , \1110 , \1111 );
mand \mul_16_12/U$1362 ( \1200 , \1112 , \1115 );
mor \mul_16_12/U$1360 ( \1201 , \1199 , \1200 );
mxor \mul_16_12/U$1356 ( \1202 , \1198 , \1201 );
mand \mul_16_12/U$1299 ( \1203 , \1035_A[3] , \979_B[2] );
mxor \mul_16_12/U$1274 ( \1204 , \1202 , \1203 );
mand \mul_16_12/U$1278 ( \1205 , \1116 , \1117 );
mand \mul_16_12/U$1277 ( \1206 , \1118 , \1121 );
mor \mul_16_12/U$1275 ( \1207 , \1205 , \1206 );
mxor \mul_16_12/U$1271 ( \1208 , \1204 , \1207 );
mand \mul_16_12/U$1207 ( \1209 , \973_A[2] , \1047_B[3] );
mxor \mul_16_12/U$1186 ( \1210 , \1208 , \1209 );
mand \mul_16_12/U$1190 ( \1211 , \1122 , \1123 );
mand \mul_16_12/U$1189 ( \1212 , \1124 , \1125 );
mor \mul_16_12/U$1187 ( \1213 , \1211 , \1212 );
mxor \mul_16_12/U$1183 ( \1214 , \1210 , \1213 );
mand \mul_16_12/U$1115 ( \1215 , \927_A[1] , \1127_B[4] );
mxor \mul_16_12/U$1098 ( \1216 , \1214 , \1215 );
mand \mul_16_12/U$1099 ( \1217 , \1126 , \1128 );
mxor \mul_16_12/U$1095 ( \1218 , \1216 , \1217 );
mbuf \mul_16_12/B[5] ( \1219_B[5] , \d[5] );
mand \mul_16_12/U$1023 ( \1220 , \891_A[0] , \1219_B[5] );
mxor \mul_16_12/U$1007 ( \1221 , \1218 , \1220 );
mbuf \mul_16_12/Z[5] ( \1222_Z[5] , \1221 );
mand \U$1/U$78 ( \1223 , \1222_Z[5] , \865 );
mbuf \add_15_12/A[5] ( \1224_A[5] , \b[5] );
mbuf \add_15_12/B[5] ( \1225_B[5] , \d[5] );
mxor \add_15_12/U$62 ( \1226 , \1224_A[5] , \1225_B[5] );
mand \add_15_12/U$66 ( \1227 , \1132_A[4] , \1133_B[4] );
mand \add_15_12/U$65 ( \1228 , \1133_B[4] , \1138 );
mand \add_15_12/U$64 ( \1229 , \1132_A[4] , \1138 );
mor \add_15_12/U$63 ( \1230 , \1227 , \1228 , \1229 );
mxor \add_15_12/U$61 ( \1231 , \1226 , \1230 );
mbuf \add_15_12/SUM[5] ( \1232_SUM[5] , \1231 );
mand \U$1/U$77 ( \1233 , \1232_SUM[5] , \863 );
mbuf \add_14_12/A[5] ( \1234_A[5] , \a[5] );
mbuf \add_14_12/B[5] ( \1235_B[5] , \c[5] );
mxor \add_14_12/U$62 ( \1236 , \1234_A[5] , \1235_B[5] );
mand \add_14_12/U$66 ( \1237 , \1142_A[4] , \1143_B[4] );
mand \add_14_12/U$65 ( \1238 , \1143_B[4] , \1148 );
mand \add_14_12/U$64 ( \1239 , \1142_A[4] , \1148 );
mor \add_14_12/U$63 ( \1240 , \1237 , \1238 , \1239 );
mxor \add_14_12/U$61 ( \1241 , \1236 , \1240 );
mbuf \add_14_12/SUM[5] ( \1242_SUM[5] , \1241 );
mand \U$1/U$76 ( \1243 , \1242_SUM[5] , \861 );
mand \U$1/U$75 ( \1244 , \d[5] , \859 );
mand \U$1/U$74 ( \1245 , \c[5] , \857 );
mand \U$1/U$73 ( \1246 , \b[5] , \855 );
mand \U$1/U$72 ( \1247 , \a[5] , \853 );
mor \U$1/U$71 ( \1248 , \1157 , \1159 , \1161 , \1163 , \1165 , \1194 , \1223 , \1233 , \1243 , \1244 , \1245 , \1246 , \1247 );
m_DC \n22[6]_g1 ( \1249 , 1'b0 , \876 );
mor \U$5/U$7 ( \1250 , \a[6] , \d[6] );
mand \U$1/U$97 ( \1251 , \1250 , \875 );
mand \U$4/U$7 ( \1252 , \b[6] , \c[6] );
mand \U$1/U$96 ( \1253 , \1252 , \873 );
mor \U$3/U$7 ( \1254 , \a[6] , \b[6] );
mand \U$1/U$95 ( \1255 , \1254 , \871 );
mxor \U$2/U$7 ( \1256 , \c[6] , \d[6] );
mand \U$1/U$94 ( \1257 , \1256 , \869 );
mbuf \mul_17_13/A[6] ( \1258_A[6] , \b[6] );
mand \mul_17_13/U$1402 ( \1259 , \1258_A[6] , \887_B[0] );
mand \mul_17_13/U$1387 ( \1260 , \1166_A[5] , \922_B[1] );
mxor \mul_17_13/U$1354 ( \1261 , \1259 , \1260 );
mand \mul_17_13/U$1358 ( \1262 , \1167 , \1168 );
mand \mul_17_13/U$1357 ( \1263 , \1169 , \1172 );
mor \mul_17_13/U$1355 ( \1264 , \1262 , \1263 );
mxor \mul_17_13/U$1351 ( \1265 , \1261 , \1264 );
mand \mul_17_13/U$1298 ( \1266 , \1086_A[4] , \968_B[2] );
mxor \mul_17_13/U$1269 ( \1267 , \1265 , \1266 );
mand \mul_17_13/U$1273 ( \1268 , \1173 , \1174 );
mand \mul_17_13/U$1272 ( \1269 , \1175 , \1178 );
mor \mul_17_13/U$1270 ( \1270 , \1268 , \1269 );
mxor \mul_17_13/U$1266 ( \1271 , \1267 , \1270 );
mand \mul_17_13/U$1206 ( \1272 , \1018_A[3] , \1030_B[3] );
mxor \mul_17_13/U$1181 ( \1273 , \1271 , \1272 );
mand \mul_17_13/U$1185 ( \1274 , \1179 , \1180 );
mand \mul_17_13/U$1184 ( \1275 , \1181 , \1184 );
mor \mul_17_13/U$1182 ( \1276 , \1274 , \1275 );
mxor \mul_17_13/U$1178 ( \1277 , \1273 , \1276 );
mand \mul_17_13/U$1114 ( \1278 , \962_A[2] , \1104_B[4] );
mxor \mul_17_13/U$1093 ( \1279 , \1277 , \1278 );
mand \mul_17_13/U$1097 ( \1280 , \1185 , \1186 );
mand \mul_17_13/U$1096 ( \1281 , \1187 , \1188 );
mor \mul_17_13/U$1094 ( \1282 , \1280 , \1281 );
mxor \mul_17_13/U$1090 ( \1283 , \1279 , \1282 );
mand \mul_17_13/U$1022 ( \1284 , \920_A[1] , \1190_B[5] );
mxor \mul_17_13/U$1005 ( \1285 , \1283 , \1284 );
mand \mul_17_13/U$1006 ( \1286 , \1189 , \1191 );
mxor \mul_17_13/U$1002 ( \1287 , \1285 , \1286 );
mbuf \mul_17_13/B[6] ( \1288_B[6] , \c[6] );
mand \mul_17_13/U$930 ( \1289 , \886_A[0] , \1288_B[6] );
mxor \mul_17_13/U$914 ( \1290 , \1287 , \1289 );
mbuf \mul_17_13/Z[6] ( \1291_Z[6] , \1290 );
mand \U$1/U$93 ( \1292 , \1291_Z[6] , \867 );
mbuf \mul_16_12/A[6] ( \1293_A[6] , \a[6] );
mand \mul_16_12/U$1402 ( \1294 , \1293_A[6] , \892_B[0] );
mand \mul_16_12/U$1387 ( \1295 , \1195_A[5] , \929_B[1] );
mxor \mul_16_12/U$1354 ( \1296 , \1294 , \1295 );
mand \mul_16_12/U$1358 ( \1297 , \1196 , \1197 );
mand \mul_16_12/U$1357 ( \1298 , \1198 , \1201 );
mor \mul_16_12/U$1355 ( \1299 , \1297 , \1298 );
mxor \mul_16_12/U$1351 ( \1300 , \1296 , \1299 );
mand \mul_16_12/U$1298 ( \1301 , \1109_A[4] , \979_B[2] );
mxor \mul_16_12/U$1269 ( \1302 , \1300 , \1301 );
mand \mul_16_12/U$1273 ( \1303 , \1202 , \1203 );
mand \mul_16_12/U$1272 ( \1304 , \1204 , \1207 );
mor \mul_16_12/U$1270 ( \1305 , \1303 , \1304 );
mxor \mul_16_12/U$1266 ( \1306 , \1302 , \1305 );
mand \mul_16_12/U$1206 ( \1307 , \1035_A[3] , \1047_B[3] );
mxor \mul_16_12/U$1181 ( \1308 , \1306 , \1307 );
mand \mul_16_12/U$1185 ( \1309 , \1208 , \1209 );
mand \mul_16_12/U$1184 ( \1310 , \1210 , \1213 );
mor \mul_16_12/U$1182 ( \1311 , \1309 , \1310 );
mxor \mul_16_12/U$1178 ( \1312 , \1308 , \1311 );
mand \mul_16_12/U$1114 ( \1313 , \973_A[2] , \1127_B[4] );
mxor \mul_16_12/U$1093 ( \1314 , \1312 , \1313 );
mand \mul_16_12/U$1097 ( \1315 , \1214 , \1215 );
mand \mul_16_12/U$1096 ( \1316 , \1216 , \1217 );
mor \mul_16_12/U$1094 ( \1317 , \1315 , \1316 );
mxor \mul_16_12/U$1090 ( \1318 , \1314 , \1317 );
mand \mul_16_12/U$1022 ( \1319 , \927_A[1] , \1219_B[5] );
mxor \mul_16_12/U$1005 ( \1320 , \1318 , \1319 );
mand \mul_16_12/U$1006 ( \1321 , \1218 , \1220 );
mxor \mul_16_12/U$1002 ( \1322 , \1320 , \1321 );
mbuf \mul_16_12/B[6] ( \1323_B[6] , \d[6] );
mand \mul_16_12/U$930 ( \1324 , \891_A[0] , \1323_B[6] );
mxor \mul_16_12/U$914 ( \1325 , \1322 , \1324 );
mbuf \mul_16_12/Z[6] ( \1326_Z[6] , \1325 );
mand \U$1/U$92 ( \1327 , \1326_Z[6] , \865 );
mbuf \add_15_12/A[6] ( \1328_A[6] , \b[6] );
mbuf \add_15_12/B[6] ( \1329_B[6] , \d[6] );
mxor \add_15_12/U$56 ( \1330 , \1328_A[6] , \1329_B[6] );
mand \add_15_12/U$60 ( \1331 , \1224_A[5] , \1225_B[5] );
mand \add_15_12/U$59 ( \1332 , \1225_B[5] , \1230 );
mand \add_15_12/U$58 ( \1333 , \1224_A[5] , \1230 );
mor \add_15_12/U$57 ( \1334 , \1331 , \1332 , \1333 );
mxor \add_15_12/U$55 ( \1335 , \1330 , \1334 );
mbuf \add_15_12/SUM[6] ( \1336_SUM[6] , \1335 );
mand \U$1/U$91 ( \1337 , \1336_SUM[6] , \863 );
mbuf \add_14_12/A[6] ( \1338_A[6] , \a[6] );
mbuf \add_14_12/B[6] ( \1339_B[6] , \c[6] );
mxor \add_14_12/U$56 ( \1340 , \1338_A[6] , \1339_B[6] );
mand \add_14_12/U$60 ( \1341 , \1234_A[5] , \1235_B[5] );
mand \add_14_12/U$59 ( \1342 , \1235_B[5] , \1240 );
mand \add_14_12/U$58 ( \1343 , \1234_A[5] , \1240 );
mor \add_14_12/U$57 ( \1344 , \1341 , \1342 , \1343 );
mxor \add_14_12/U$55 ( \1345 , \1340 , \1344 );
mbuf \add_14_12/SUM[6] ( \1346_SUM[6] , \1345 );
mand \U$1/U$90 ( \1347 , \1346_SUM[6] , \861 );
mand \U$1/U$89 ( \1348 , \d[6] , \859 );
mand \U$1/U$88 ( \1349 , \c[6] , \857 );
mand \U$1/U$87 ( \1350 , \b[6] , \855 );
mand \U$1/U$86 ( \1351 , \a[6] , \853 );
mor \U$1/U$85 ( \1352 , \1249 , \1251 , \1253 , \1255 , \1257 , \1292 , \1327 , \1337 , \1347 , \1348 , \1349 , \1350 , \1351 );
m_DC \n22[7]_g1 ( \1353 , 1'b0 , \876 );
mor \U$5/U$8 ( \1354 , \a[7] , \d[7] );
mand \U$1/U$111 ( \1355 , \1354 , \875 );
mand \U$4/U$8 ( \1356 , \b[7] , \c[7] );
mand \U$1/U$110 ( \1357 , \1356 , \873 );
mor \U$3/U$8 ( \1358 , \a[7] , \b[7] );
mand \U$1/U$109 ( \1359 , \1358 , \871 );
mxor \U$2/U$8 ( \1360 , \c[7] , \d[7] );
mand \U$1/U$108 ( \1361 , \1360 , \869 );
mbuf \mul_17_13/A[7] ( \1362_A[7] , \b[7] );
mand \mul_17_13/U$1401 ( \1363 , \1362_A[7] , \887_B[0] );
mand \mul_17_13/U$1386 ( \1364 , \1258_A[6] , \922_B[1] );
mxor \mul_17_13/U$1349 ( \1365 , \1363 , \1364 );
mand \mul_17_13/U$1353 ( \1366 , \1259 , \1260 );
mand \mul_17_13/U$1352 ( \1367 , \1261 , \1264 );
mor \mul_17_13/U$1350 ( \1368 , \1366 , \1367 );
mxor \mul_17_13/U$1346 ( \1369 , \1365 , \1368 );
mand \mul_17_13/U$1297 ( \1370 , \1166_A[5] , \968_B[2] );
mxor \mul_17_13/U$1264 ( \1371 , \1369 , \1370 );
mand \mul_17_13/U$1268 ( \1372 , \1265 , \1266 );
mand \mul_17_13/U$1267 ( \1373 , \1267 , \1270 );
mor \mul_17_13/U$1265 ( \1374 , \1372 , \1373 );
mxor \mul_17_13/U$1261 ( \1375 , \1371 , \1374 );
mand \mul_17_13/U$1205 ( \1376 , \1086_A[4] , \1030_B[3] );
mxor \mul_17_13/U$1176 ( \1377 , \1375 , \1376 );
mand \mul_17_13/U$1180 ( \1378 , \1271 , \1272 );
mand \mul_17_13/U$1179 ( \1379 , \1273 , \1276 );
mor \mul_17_13/U$1177 ( \1380 , \1378 , \1379 );
mxor \mul_17_13/U$1173 ( \1381 , \1377 , \1380 );
mand \mul_17_13/U$1113 ( \1382 , \1018_A[3] , \1104_B[4] );
mxor \mul_17_13/U$1088 ( \1383 , \1381 , \1382 );
mand \mul_17_13/U$1092 ( \1384 , \1277 , \1278 );
mand \mul_17_13/U$1091 ( \1385 , \1279 , \1282 );
mor \mul_17_13/U$1089 ( \1386 , \1384 , \1385 );
mxor \mul_17_13/U$1085 ( \1387 , \1383 , \1386 );
mand \mul_17_13/U$1021 ( \1388 , \962_A[2] , \1190_B[5] );
mxor \mul_17_13/U$1000 ( \1389 , \1387 , \1388 );
mand \mul_17_13/U$1004 ( \1390 , \1283 , \1284 );
mand \mul_17_13/U$1003 ( \1391 , \1285 , \1286 );
mor \mul_17_13/U$1001 ( \1392 , \1390 , \1391 );
mxor \mul_17_13/U$997 ( \1393 , \1389 , \1392 );
mand \mul_17_13/U$929 ( \1394 , \920_A[1] , \1288_B[6] );
mxor \mul_17_13/U$912 ( \1395 , \1393 , \1394 );
mand \mul_17_13/U$913 ( \1396 , \1287 , \1289 );
mxor \mul_17_13/U$909 ( \1397 , \1395 , \1396 );
mbuf \mul_17_13/B[7] ( \1398_B[7] , \c[7] );
mand \mul_17_13/U$837 ( \1399 , \886_A[0] , \1398_B[7] );
mxor \mul_17_13/U$821 ( \1400 , \1397 , \1399 );
mbuf \mul_17_13/Z[7] ( \1401_Z[7] , \1400 );
mand \U$1/U$107 ( \1402 , \1401_Z[7] , \867 );
mbuf \mul_16_12/A[7] ( \1403_A[7] , \a[7] );
mand \mul_16_12/U$1401 ( \1404 , \1403_A[7] , \892_B[0] );
mand \mul_16_12/U$1386 ( \1405 , \1293_A[6] , \929_B[1] );
mxor \mul_16_12/U$1349 ( \1406 , \1404 , \1405 );
mand \mul_16_12/U$1353 ( \1407 , \1294 , \1295 );
mand \mul_16_12/U$1352 ( \1408 , \1296 , \1299 );
mor \mul_16_12/U$1350 ( \1409 , \1407 , \1408 );
mxor \mul_16_12/U$1346 ( \1410 , \1406 , \1409 );
mand \mul_16_12/U$1297 ( \1411 , \1195_A[5] , \979_B[2] );
mxor \mul_16_12/U$1264 ( \1412 , \1410 , \1411 );
mand \mul_16_12/U$1268 ( \1413 , \1300 , \1301 );
mand \mul_16_12/U$1267 ( \1414 , \1302 , \1305 );
mor \mul_16_12/U$1265 ( \1415 , \1413 , \1414 );
mxor \mul_16_12/U$1261 ( \1416 , \1412 , \1415 );
mand \mul_16_12/U$1205 ( \1417 , \1109_A[4] , \1047_B[3] );
mxor \mul_16_12/U$1176 ( \1418 , \1416 , \1417 );
mand \mul_16_12/U$1180 ( \1419 , \1306 , \1307 );
mand \mul_16_12/U$1179 ( \1420 , \1308 , \1311 );
mor \mul_16_12/U$1177 ( \1421 , \1419 , \1420 );
mxor \mul_16_12/U$1173 ( \1422 , \1418 , \1421 );
mand \mul_16_12/U$1113 ( \1423 , \1035_A[3] , \1127_B[4] );
mxor \mul_16_12/U$1088 ( \1424 , \1422 , \1423 );
mand \mul_16_12/U$1092 ( \1425 , \1312 , \1313 );
mand \mul_16_12/U$1091 ( \1426 , \1314 , \1317 );
mor \mul_16_12/U$1089 ( \1427 , \1425 , \1426 );
mxor \mul_16_12/U$1085 ( \1428 , \1424 , \1427 );
mand \mul_16_12/U$1021 ( \1429 , \973_A[2] , \1219_B[5] );
mxor \mul_16_12/U$1000 ( \1430 , \1428 , \1429 );
mand \mul_16_12/U$1004 ( \1431 , \1318 , \1319 );
mand \mul_16_12/U$1003 ( \1432 , \1320 , \1321 );
mor \mul_16_12/U$1001 ( \1433 , \1431 , \1432 );
mxor \mul_16_12/U$997 ( \1434 , \1430 , \1433 );
mand \mul_16_12/U$929 ( \1435 , \927_A[1] , \1323_B[6] );
mxor \mul_16_12/U$912 ( \1436 , \1434 , \1435 );
mand \mul_16_12/U$913 ( \1437 , \1322 , \1324 );
mxor \mul_16_12/U$909 ( \1438 , \1436 , \1437 );
mbuf \mul_16_12/B[7] ( \1439_B[7] , \d[7] );
mand \mul_16_12/U$837 ( \1440 , \891_A[0] , \1439_B[7] );
mxor \mul_16_12/U$821 ( \1441 , \1438 , \1440 );
mbuf \mul_16_12/Z[7] ( \1442_Z[7] , \1441 );
mand \U$1/U$106 ( \1443 , \1442_Z[7] , \865 );
mbuf \add_15_12/A[7] ( \1444_A[7] , \b[7] );
mbuf \add_15_12/B[7] ( \1445_B[7] , \d[7] );
mxor \add_15_12/U$50 ( \1446 , \1444_A[7] , \1445_B[7] );
mand \add_15_12/U$54 ( \1447 , \1328_A[6] , \1329_B[6] );
mand \add_15_12/U$53 ( \1448 , \1329_B[6] , \1334 );
mand \add_15_12/U$52 ( \1449 , \1328_A[6] , \1334 );
mor \add_15_12/U$51 ( \1450 , \1447 , \1448 , \1449 );
mxor \add_15_12/U$49 ( \1451 , \1446 , \1450 );
mbuf \add_15_12/SUM[7] ( \1452_SUM[7] , \1451 );
mand \U$1/U$105 ( \1453 , \1452_SUM[7] , \863 );
mbuf \add_14_12/A[7] ( \1454_A[7] , \a[7] );
mbuf \add_14_12/B[7] ( \1455_B[7] , \c[7] );
mxor \add_14_12/U$50 ( \1456 , \1454_A[7] , \1455_B[7] );
mand \add_14_12/U$54 ( \1457 , \1338_A[6] , \1339_B[6] );
mand \add_14_12/U$53 ( \1458 , \1339_B[6] , \1344 );
mand \add_14_12/U$52 ( \1459 , \1338_A[6] , \1344 );
mor \add_14_12/U$51 ( \1460 , \1457 , \1458 , \1459 );
mxor \add_14_12/U$49 ( \1461 , \1456 , \1460 );
mbuf \add_14_12/SUM[7] ( \1462_SUM[7] , \1461 );
mand \U$1/U$104 ( \1463 , \1462_SUM[7] , \861 );
mand \U$1/U$103 ( \1464 , \d[7] , \859 );
mand \U$1/U$102 ( \1465 , \c[7] , \857 );
mand \U$1/U$101 ( \1466 , \b[7] , \855 );
mand \U$1/U$100 ( \1467 , \a[7] , \853 );
mor \U$1/U$99 ( \1468 , \1353 , \1355 , \1357 , \1359 , \1361 , \1402 , \1443 , \1453 , \1463 , \1464 , \1465 , \1466 , \1467 );
m_DC \n22[8]_g1 ( \1469 , 1'b0 , \876 );
mor \U$5/U$9 ( \1470 , \a[8] , \d[8] );
mand \U$1/U$125 ( \1471 , \1470 , \875 );
mand \U$4/U$9 ( \1472 , \b[8] , \c[8] );
mand \U$1/U$124 ( \1473 , \1472 , \873 );
mor \U$3/U$9 ( \1474 , \a[8] , \b[8] );
mand \U$1/U$123 ( \1475 , \1474 , \871 );
mxor \U$2/U$9 ( \1476 , \c[8] , \d[8] );
mand \U$1/U$122 ( \1477 , \1476 , \869 );
mbuf \mul_17_13/A[8] ( \1478_A[8] , \b[8] );
mand \mul_17_13/U$1400 ( \1479 , \1478_A[8] , \887_B[0] );
mand \mul_17_13/U$1385 ( \1480 , \1362_A[7] , \922_B[1] );
mxor \mul_17_13/U$1344 ( \1481 , \1479 , \1480 );
mand \mul_17_13/U$1348 ( \1482 , \1363 , \1364 );
mand \mul_17_13/U$1347 ( \1483 , \1365 , \1368 );
mor \mul_17_13/U$1345 ( \1484 , \1482 , \1483 );
mxor \mul_17_13/U$1341 ( \1485 , \1481 , \1484 );
mand \mul_17_13/U$1296 ( \1486 , \1258_A[6] , \968_B[2] );
mxor \mul_17_13/U$1259 ( \1487 , \1485 , \1486 );
mand \mul_17_13/U$1263 ( \1488 , \1369 , \1370 );
mand \mul_17_13/U$1262 ( \1489 , \1371 , \1374 );
mor \mul_17_13/U$1260 ( \1490 , \1488 , \1489 );
mxor \mul_17_13/U$1256 ( \1491 , \1487 , \1490 );
mand \mul_17_13/U$1204 ( \1492 , \1166_A[5] , \1030_B[3] );
mxor \mul_17_13/U$1171 ( \1493 , \1491 , \1492 );
mand \mul_17_13/U$1175 ( \1494 , \1375 , \1376 );
mand \mul_17_13/U$1174 ( \1495 , \1377 , \1380 );
mor \mul_17_13/U$1172 ( \1496 , \1494 , \1495 );
mxor \mul_17_13/U$1168 ( \1497 , \1493 , \1496 );
mand \mul_17_13/U$1112 ( \1498 , \1086_A[4] , \1104_B[4] );
mxor \mul_17_13/U$1083 ( \1499 , \1497 , \1498 );
mand \mul_17_13/U$1087 ( \1500 , \1381 , \1382 );
mand \mul_17_13/U$1086 ( \1501 , \1383 , \1386 );
mor \mul_17_13/U$1084 ( \1502 , \1500 , \1501 );
mxor \mul_17_13/U$1080 ( \1503 , \1499 , \1502 );
mand \mul_17_13/U$1020 ( \1504 , \1018_A[3] , \1190_B[5] );
mxor \mul_17_13/U$995 ( \1505 , \1503 , \1504 );
mand \mul_17_13/U$999 ( \1506 , \1387 , \1388 );
mand \mul_17_13/U$998 ( \1507 , \1389 , \1392 );
mor \mul_17_13/U$996 ( \1508 , \1506 , \1507 );
mxor \mul_17_13/U$992 ( \1509 , \1505 , \1508 );
mand \mul_17_13/U$928 ( \1510 , \962_A[2] , \1288_B[6] );
mxor \mul_17_13/U$907 ( \1511 , \1509 , \1510 );
mand \mul_17_13/U$911 ( \1512 , \1393 , \1394 );
mand \mul_17_13/U$910 ( \1513 , \1395 , \1396 );
mor \mul_17_13/U$908 ( \1514 , \1512 , \1513 );
mxor \mul_17_13/U$904 ( \1515 , \1511 , \1514 );
mand \mul_17_13/U$836 ( \1516 , \920_A[1] , \1398_B[7] );
mxor \mul_17_13/U$819 ( \1517 , \1515 , \1516 );
mand \mul_17_13/U$820 ( \1518 , \1397 , \1399 );
mxor \mul_17_13/U$816 ( \1519 , \1517 , \1518 );
mbuf \mul_17_13/B[8] ( \1520_B[8] , \c[8] );
mand \mul_17_13/U$744 ( \1521 , \886_A[0] , \1520_B[8] );
mxor \mul_17_13/U$728 ( \1522 , \1519 , \1521 );
mbuf \mul_17_13/Z[8] ( \1523_Z[8] , \1522 );
mand \U$1/U$121 ( \1524 , \1523_Z[8] , \867 );
mbuf \mul_16_12/A[8] ( \1525_A[8] , \a[8] );
mand \mul_16_12/U$1400 ( \1526 , \1525_A[8] , \892_B[0] );
mand \mul_16_12/U$1385 ( \1527 , \1403_A[7] , \929_B[1] );
mxor \mul_16_12/U$1344 ( \1528 , \1526 , \1527 );
mand \mul_16_12/U$1348 ( \1529 , \1404 , \1405 );
mand \mul_16_12/U$1347 ( \1530 , \1406 , \1409 );
mor \mul_16_12/U$1345 ( \1531 , \1529 , \1530 );
mxor \mul_16_12/U$1341 ( \1532 , \1528 , \1531 );
mand \mul_16_12/U$1296 ( \1533 , \1293_A[6] , \979_B[2] );
mxor \mul_16_12/U$1259 ( \1534 , \1532 , \1533 );
mand \mul_16_12/U$1263 ( \1535 , \1410 , \1411 );
mand \mul_16_12/U$1262 ( \1536 , \1412 , \1415 );
mor \mul_16_12/U$1260 ( \1537 , \1535 , \1536 );
mxor \mul_16_12/U$1256 ( \1538 , \1534 , \1537 );
mand \mul_16_12/U$1204 ( \1539 , \1195_A[5] , \1047_B[3] );
mxor \mul_16_12/U$1171 ( \1540 , \1538 , \1539 );
mand \mul_16_12/U$1175 ( \1541 , \1416 , \1417 );
mand \mul_16_12/U$1174 ( \1542 , \1418 , \1421 );
mor \mul_16_12/U$1172 ( \1543 , \1541 , \1542 );
mxor \mul_16_12/U$1168 ( \1544 , \1540 , \1543 );
mand \mul_16_12/U$1112 ( \1545 , \1109_A[4] , \1127_B[4] );
mxor \mul_16_12/U$1083 ( \1546 , \1544 , \1545 );
mand \mul_16_12/U$1087 ( \1547 , \1422 , \1423 );
mand \mul_16_12/U$1086 ( \1548 , \1424 , \1427 );
mor \mul_16_12/U$1084 ( \1549 , \1547 , \1548 );
mxor \mul_16_12/U$1080 ( \1550 , \1546 , \1549 );
mand \mul_16_12/U$1020 ( \1551 , \1035_A[3] , \1219_B[5] );
mxor \mul_16_12/U$995 ( \1552 , \1550 , \1551 );
mand \mul_16_12/U$999 ( \1553 , \1428 , \1429 );
mand \mul_16_12/U$998 ( \1554 , \1430 , \1433 );
mor \mul_16_12/U$996 ( \1555 , \1553 , \1554 );
mxor \mul_16_12/U$992 ( \1556 , \1552 , \1555 );
mand \mul_16_12/U$928 ( \1557 , \973_A[2] , \1323_B[6] );
mxor \mul_16_12/U$907 ( \1558 , \1556 , \1557 );
mand \mul_16_12/U$911 ( \1559 , \1434 , \1435 );
mand \mul_16_12/U$910 ( \1560 , \1436 , \1437 );
mor \mul_16_12/U$908 ( \1561 , \1559 , \1560 );
mxor \mul_16_12/U$904 ( \1562 , \1558 , \1561 );
mand \mul_16_12/U$836 ( \1563 , \927_A[1] , \1439_B[7] );
mxor \mul_16_12/U$819 ( \1564 , \1562 , \1563 );
mand \mul_16_12/U$820 ( \1565 , \1438 , \1440 );
mxor \mul_16_12/U$816 ( \1566 , \1564 , \1565 );
mbuf \mul_16_12/B[8] ( \1567_B[8] , \d[8] );
mand \mul_16_12/U$744 ( \1568 , \891_A[0] , \1567_B[8] );
mxor \mul_16_12/U$728 ( \1569 , \1566 , \1568 );
mbuf \mul_16_12/Z[8] ( \1570_Z[8] , \1569 );
mand \U$1/U$120 ( \1571 , \1570_Z[8] , \865 );
mbuf \add_15_12/A[8] ( \1572_A[8] , \b[8] );
mbuf \add_15_12/B[8] ( \1573_B[8] , \d[8] );
mxor \add_15_12/U$44 ( \1574 , \1572_A[8] , \1573_B[8] );
mand \add_15_12/U$48 ( \1575 , \1444_A[7] , \1445_B[7] );
mand \add_15_12/U$47 ( \1576 , \1445_B[7] , \1450 );
mand \add_15_12/U$46 ( \1577 , \1444_A[7] , \1450 );
mor \add_15_12/U$45 ( \1578 , \1575 , \1576 , \1577 );
mxor \add_15_12/U$43 ( \1579 , \1574 , \1578 );
mbuf \add_15_12/SUM[8] ( \1580_SUM[8] , \1579 );
mand \U$1/U$119 ( \1581 , \1580_SUM[8] , \863 );
mbuf \add_14_12/A[8] ( \1582_A[8] , \a[8] );
mbuf \add_14_12/B[8] ( \1583_B[8] , \c[8] );
mxor \add_14_12/U$44 ( \1584 , \1582_A[8] , \1583_B[8] );
mand \add_14_12/U$48 ( \1585 , \1454_A[7] , \1455_B[7] );
mand \add_14_12/U$47 ( \1586 , \1455_B[7] , \1460 );
mand \add_14_12/U$46 ( \1587 , \1454_A[7] , \1460 );
mor \add_14_12/U$45 ( \1588 , \1585 , \1586 , \1587 );
mxor \add_14_12/U$43 ( \1589 , \1584 , \1588 );
mbuf \add_14_12/SUM[8] ( \1590_SUM[8] , \1589 );
mand \U$1/U$118 ( \1591 , \1590_SUM[8] , \861 );
mand \U$1/U$117 ( \1592 , \d[8] , \859 );
mand \U$1/U$116 ( \1593 , \c[8] , \857 );
mand \U$1/U$115 ( \1594 , \b[8] , \855 );
mand \U$1/U$114 ( \1595 , \a[8] , \853 );
mor \U$1/U$113 ( \1596 , \1469 , \1471 , \1473 , \1475 , \1477 , \1524 , \1571 , \1581 , \1591 , \1592 , \1593 , \1594 , \1595 );
m_DC \n22[9]_g1 ( \1597 , 1'b0 , \876 );
mor \U$5/U$10 ( \1598 , \a[9] , \d[9] );
mand \U$1/U$139 ( \1599 , \1598 , \875 );
mand \U$4/U$10 ( \1600 , \b[9] , \c[9] );
mand \U$1/U$138 ( \1601 , \1600 , \873 );
mor \U$3/U$10 ( \1602 , \a[9] , \b[9] );
mand \U$1/U$137 ( \1603 , \1602 , \871 );
mxor \U$2/U$10 ( \1604 , \c[9] , \d[9] );
mand \U$1/U$136 ( \1605 , \1604 , \869 );
mbuf \mul_17_13/A[9] ( \1606_A[9] , \b[9] );
mand \mul_17_13/U$1399 ( \1607 , \1606_A[9] , \887_B[0] );
mand \mul_17_13/U$1384 ( \1608 , \1478_A[8] , \922_B[1] );
mxor \mul_17_13/U$1339 ( \1609 , \1607 , \1608 );
mand \mul_17_13/U$1343 ( \1610 , \1479 , \1480 );
mand \mul_17_13/U$1342 ( \1611 , \1481 , \1484 );
mor \mul_17_13/U$1340 ( \1612 , \1610 , \1611 );
mxor \mul_17_13/U$1336 ( \1613 , \1609 , \1612 );
mand \mul_17_13/U$1295 ( \1614 , \1362_A[7] , \968_B[2] );
mxor \mul_17_13/U$1254 ( \1615 , \1613 , \1614 );
mand \mul_17_13/U$1258 ( \1616 , \1485 , \1486 );
mand \mul_17_13/U$1257 ( \1617 , \1487 , \1490 );
mor \mul_17_13/U$1255 ( \1618 , \1616 , \1617 );
mxor \mul_17_13/U$1251 ( \1619 , \1615 , \1618 );
mand \mul_17_13/U$1203 ( \1620 , \1258_A[6] , \1030_B[3] );
mxor \mul_17_13/U$1166 ( \1621 , \1619 , \1620 );
mand \mul_17_13/U$1170 ( \1622 , \1491 , \1492 );
mand \mul_17_13/U$1169 ( \1623 , \1493 , \1496 );
mor \mul_17_13/U$1167 ( \1624 , \1622 , \1623 );
mxor \mul_17_13/U$1163 ( \1625 , \1621 , \1624 );
mand \mul_17_13/U$1111 ( \1626 , \1166_A[5] , \1104_B[4] );
mxor \mul_17_13/U$1078 ( \1627 , \1625 , \1626 );
mand \mul_17_13/U$1082 ( \1628 , \1497 , \1498 );
mand \mul_17_13/U$1081 ( \1629 , \1499 , \1502 );
mor \mul_17_13/U$1079 ( \1630 , \1628 , \1629 );
mxor \mul_17_13/U$1075 ( \1631 , \1627 , \1630 );
mand \mul_17_13/U$1019 ( \1632 , \1086_A[4] , \1190_B[5] );
mxor \mul_17_13/U$990 ( \1633 , \1631 , \1632 );
mand \mul_17_13/U$994 ( \1634 , \1503 , \1504 );
mand \mul_17_13/U$993 ( \1635 , \1505 , \1508 );
mor \mul_17_13/U$991 ( \1636 , \1634 , \1635 );
mxor \mul_17_13/U$987 ( \1637 , \1633 , \1636 );
mand \mul_17_13/U$927 ( \1638 , \1018_A[3] , \1288_B[6] );
mxor \mul_17_13/U$902 ( \1639 , \1637 , \1638 );
mand \mul_17_13/U$906 ( \1640 , \1509 , \1510 );
mand \mul_17_13/U$905 ( \1641 , \1511 , \1514 );
mor \mul_17_13/U$903 ( \1642 , \1640 , \1641 );
mxor \mul_17_13/U$899 ( \1643 , \1639 , \1642 );
mand \mul_17_13/U$835 ( \1644 , \962_A[2] , \1398_B[7] );
mxor \mul_17_13/U$814 ( \1645 , \1643 , \1644 );
mand \mul_17_13/U$818 ( \1646 , \1515 , \1516 );
mand \mul_17_13/U$817 ( \1647 , \1517 , \1518 );
mor \mul_17_13/U$815 ( \1648 , \1646 , \1647 );
mxor \mul_17_13/U$811 ( \1649 , \1645 , \1648 );
mand \mul_17_13/U$743 ( \1650 , \920_A[1] , \1520_B[8] );
mxor \mul_17_13/U$726 ( \1651 , \1649 , \1650 );
mand \mul_17_13/U$727 ( \1652 , \1519 , \1521 );
mxor \mul_17_13/U$723 ( \1653 , \1651 , \1652 );
mbuf \mul_17_13/B[9] ( \1654_B[9] , \c[9] );
mand \mul_17_13/U$651 ( \1655 , \886_A[0] , \1654_B[9] );
mxor \mul_17_13/U$635 ( \1656 , \1653 , \1655 );
mbuf \mul_17_13/Z[9] ( \1657_Z[9] , \1656 );
mand \U$1/U$135 ( \1658 , \1657_Z[9] , \867 );
mbuf \mul_16_12/A[9] ( \1659_A[9] , \a[9] );
mand \mul_16_12/U$1399 ( \1660 , \1659_A[9] , \892_B[0] );
mand \mul_16_12/U$1384 ( \1661 , \1525_A[8] , \929_B[1] );
mxor \mul_16_12/U$1339 ( \1662 , \1660 , \1661 );
mand \mul_16_12/U$1343 ( \1663 , \1526 , \1527 );
mand \mul_16_12/U$1342 ( \1664 , \1528 , \1531 );
mor \mul_16_12/U$1340 ( \1665 , \1663 , \1664 );
mxor \mul_16_12/U$1336 ( \1666 , \1662 , \1665 );
mand \mul_16_12/U$1295 ( \1667 , \1403_A[7] , \979_B[2] );
mxor \mul_16_12/U$1254 ( \1668 , \1666 , \1667 );
mand \mul_16_12/U$1258 ( \1669 , \1532 , \1533 );
mand \mul_16_12/U$1257 ( \1670 , \1534 , \1537 );
mor \mul_16_12/U$1255 ( \1671 , \1669 , \1670 );
mxor \mul_16_12/U$1251 ( \1672 , \1668 , \1671 );
mand \mul_16_12/U$1203 ( \1673 , \1293_A[6] , \1047_B[3] );
mxor \mul_16_12/U$1166 ( \1674 , \1672 , \1673 );
mand \mul_16_12/U$1170 ( \1675 , \1538 , \1539 );
mand \mul_16_12/U$1169 ( \1676 , \1540 , \1543 );
mor \mul_16_12/U$1167 ( \1677 , \1675 , \1676 );
mxor \mul_16_12/U$1163 ( \1678 , \1674 , \1677 );
mand \mul_16_12/U$1111 ( \1679 , \1195_A[5] , \1127_B[4] );
mxor \mul_16_12/U$1078 ( \1680 , \1678 , \1679 );
mand \mul_16_12/U$1082 ( \1681 , \1544 , \1545 );
mand \mul_16_12/U$1081 ( \1682 , \1546 , \1549 );
mor \mul_16_12/U$1079 ( \1683 , \1681 , \1682 );
mxor \mul_16_12/U$1075 ( \1684 , \1680 , \1683 );
mand \mul_16_12/U$1019 ( \1685 , \1109_A[4] , \1219_B[5] );
mxor \mul_16_12/U$990 ( \1686 , \1684 , \1685 );
mand \mul_16_12/U$994 ( \1687 , \1550 , \1551 );
mand \mul_16_12/U$993 ( \1688 , \1552 , \1555 );
mor \mul_16_12/U$991 ( \1689 , \1687 , \1688 );
mxor \mul_16_12/U$987 ( \1690 , \1686 , \1689 );
mand \mul_16_12/U$927 ( \1691 , \1035_A[3] , \1323_B[6] );
mxor \mul_16_12/U$902 ( \1692 , \1690 , \1691 );
mand \mul_16_12/U$906 ( \1693 , \1556 , \1557 );
mand \mul_16_12/U$905 ( \1694 , \1558 , \1561 );
mor \mul_16_12/U$903 ( \1695 , \1693 , \1694 );
mxor \mul_16_12/U$899 ( \1696 , \1692 , \1695 );
mand \mul_16_12/U$835 ( \1697 , \973_A[2] , \1439_B[7] );
mxor \mul_16_12/U$814 ( \1698 , \1696 , \1697 );
mand \mul_16_12/U$818 ( \1699 , \1562 , \1563 );
mand \mul_16_12/U$817 ( \1700 , \1564 , \1565 );
mor \mul_16_12/U$815 ( \1701 , \1699 , \1700 );
mxor \mul_16_12/U$811 ( \1702 , \1698 , \1701 );
mand \mul_16_12/U$743 ( \1703 , \927_A[1] , \1567_B[8] );
mxor \mul_16_12/U$726 ( \1704 , \1702 , \1703 );
mand \mul_16_12/U$727 ( \1705 , \1566 , \1568 );
mxor \mul_16_12/U$723 ( \1706 , \1704 , \1705 );
mbuf \mul_16_12/B[9] ( \1707_B[9] , \d[9] );
mand \mul_16_12/U$651 ( \1708 , \891_A[0] , \1707_B[9] );
mxor \mul_16_12/U$635 ( \1709 , \1706 , \1708 );
mbuf \mul_16_12/Z[9] ( \1710_Z[9] , \1709 );
mand \U$1/U$134 ( \1711 , \1710_Z[9] , \865 );
mbuf \add_15_12/A[9] ( \1712_A[9] , \b[9] );
mbuf \add_15_12/B[9] ( \1713_B[9] , \d[9] );
mxor \add_15_12/U$38 ( \1714 , \1712_A[9] , \1713_B[9] );
mand \add_15_12/U$42 ( \1715 , \1572_A[8] , \1573_B[8] );
mand \add_15_12/U$41 ( \1716 , \1573_B[8] , \1578 );
mand \add_15_12/U$40 ( \1717 , \1572_A[8] , \1578 );
mor \add_15_12/U$39 ( \1718 , \1715 , \1716 , \1717 );
mxor \add_15_12/U$37 ( \1719 , \1714 , \1718 );
mbuf \add_15_12/SUM[9] ( \1720_SUM[9] , \1719 );
mand \U$1/U$133 ( \1721 , \1720_SUM[9] , \863 );
mbuf \add_14_12/A[9] ( \1722_A[9] , \a[9] );
mbuf \add_14_12/B[9] ( \1723_B[9] , \c[9] );
mxor \add_14_12/U$38 ( \1724 , \1722_A[9] , \1723_B[9] );
mand \add_14_12/U$42 ( \1725 , \1582_A[8] , \1583_B[8] );
mand \add_14_12/U$41 ( \1726 , \1583_B[8] , \1588 );
mand \add_14_12/U$40 ( \1727 , \1582_A[8] , \1588 );
mor \add_14_12/U$39 ( \1728 , \1725 , \1726 , \1727 );
mxor \add_14_12/U$37 ( \1729 , \1724 , \1728 );
mbuf \add_14_12/SUM[9] ( \1730_SUM[9] , \1729 );
mand \U$1/U$132 ( \1731 , \1730_SUM[9] , \861 );
mand \U$1/U$131 ( \1732 , \d[9] , \859 );
mand \U$1/U$130 ( \1733 , \c[9] , \857 );
mand \U$1/U$129 ( \1734 , \b[9] , \855 );
mand \U$1/U$128 ( \1735 , \a[9] , \853 );
mor \U$1/U$127 ( \1736 , \1597 , \1599 , \1601 , \1603 , \1605 , \1658 , \1711 , \1721 , \1731 , \1732 , \1733 , \1734 , \1735 );
m_DC \n22[10]_g1 ( \1737 , 1'b0 , \876 );
mor \U$5/U$11 ( \1738 , \a[10] , \d[10] );
mand \U$1/U$153 ( \1739 , \1738 , \875 );
mand \U$4/U$11 ( \1740 , \b[10] , \c[10] );
mand \U$1/U$152 ( \1741 , \1740 , \873 );
mor \U$3/U$11 ( \1742 , \a[10] , \b[10] );
mand \U$1/U$151 ( \1743 , \1742 , \871 );
mxor \U$2/U$11 ( \1744 , \c[10] , \d[10] );
mand \U$1/U$150 ( \1745 , \1744 , \869 );
mbuf \mul_17_13/A[10] ( \1746_A[10] , \b[10] );
mand \mul_17_13/U$1398 ( \1747 , \1746_A[10] , \887_B[0] );
mand \mul_17_13/U$1383 ( \1748 , \1606_A[9] , \922_B[1] );
mxor \mul_17_13/U$1334 ( \1749 , \1747 , \1748 );
mand \mul_17_13/U$1338 ( \1750 , \1607 , \1608 );
mand \mul_17_13/U$1337 ( \1751 , \1609 , \1612 );
mor \mul_17_13/U$1335 ( \1752 , \1750 , \1751 );
mxor \mul_17_13/U$1331 ( \1753 , \1749 , \1752 );
mand \mul_17_13/U$1294 ( \1754 , \1478_A[8] , \968_B[2] );
mxor \mul_17_13/U$1249 ( \1755 , \1753 , \1754 );
mand \mul_17_13/U$1253 ( \1756 , \1613 , \1614 );
mand \mul_17_13/U$1252 ( \1757 , \1615 , \1618 );
mor \mul_17_13/U$1250 ( \1758 , \1756 , \1757 );
mxor \mul_17_13/U$1246 ( \1759 , \1755 , \1758 );
mand \mul_17_13/U$1202 ( \1760 , \1362_A[7] , \1030_B[3] );
mxor \mul_17_13/U$1161 ( \1761 , \1759 , \1760 );
mand \mul_17_13/U$1165 ( \1762 , \1619 , \1620 );
mand \mul_17_13/U$1164 ( \1763 , \1621 , \1624 );
mor \mul_17_13/U$1162 ( \1764 , \1762 , \1763 );
mxor \mul_17_13/U$1158 ( \1765 , \1761 , \1764 );
mand \mul_17_13/U$1110 ( \1766 , \1258_A[6] , \1104_B[4] );
mxor \mul_17_13/U$1073 ( \1767 , \1765 , \1766 );
mand \mul_17_13/U$1077 ( \1768 , \1625 , \1626 );
mand \mul_17_13/U$1076 ( \1769 , \1627 , \1630 );
mor \mul_17_13/U$1074 ( \1770 , \1768 , \1769 );
mxor \mul_17_13/U$1070 ( \1771 , \1767 , \1770 );
mand \mul_17_13/U$1018 ( \1772 , \1166_A[5] , \1190_B[5] );
mxor \mul_17_13/U$985 ( \1773 , \1771 , \1772 );
mand \mul_17_13/U$989 ( \1774 , \1631 , \1632 );
mand \mul_17_13/U$988 ( \1775 , \1633 , \1636 );
mor \mul_17_13/U$986 ( \1776 , \1774 , \1775 );
mxor \mul_17_13/U$982 ( \1777 , \1773 , \1776 );
mand \mul_17_13/U$926 ( \1778 , \1086_A[4] , \1288_B[6] );
mxor \mul_17_13/U$897 ( \1779 , \1777 , \1778 );
mand \mul_17_13/U$901 ( \1780 , \1637 , \1638 );
mand \mul_17_13/U$900 ( \1781 , \1639 , \1642 );
mor \mul_17_13/U$898 ( \1782 , \1780 , \1781 );
mxor \mul_17_13/U$894 ( \1783 , \1779 , \1782 );
mand \mul_17_13/U$834 ( \1784 , \1018_A[3] , \1398_B[7] );
mxor \mul_17_13/U$809 ( \1785 , \1783 , \1784 );
mand \mul_17_13/U$813 ( \1786 , \1643 , \1644 );
mand \mul_17_13/U$812 ( \1787 , \1645 , \1648 );
mor \mul_17_13/U$810 ( \1788 , \1786 , \1787 );
mxor \mul_17_13/U$806 ( \1789 , \1785 , \1788 );
mand \mul_17_13/U$742 ( \1790 , \962_A[2] , \1520_B[8] );
mxor \mul_17_13/U$721 ( \1791 , \1789 , \1790 );
mand \mul_17_13/U$725 ( \1792 , \1649 , \1650 );
mand \mul_17_13/U$724 ( \1793 , \1651 , \1652 );
mor \mul_17_13/U$722 ( \1794 , \1792 , \1793 );
mxor \mul_17_13/U$718 ( \1795 , \1791 , \1794 );
mand \mul_17_13/U$650 ( \1796 , \920_A[1] , \1654_B[9] );
mxor \mul_17_13/U$633 ( \1797 , \1795 , \1796 );
mand \mul_17_13/U$634 ( \1798 , \1653 , \1655 );
mxor \mul_17_13/U$630 ( \1799 , \1797 , \1798 );
mbuf \mul_17_13/B[10] ( \1800_B[10] , \c[10] );
mand \mul_17_13/U$558 ( \1801 , \886_A[0] , \1800_B[10] );
mxor \mul_17_13/U$542 ( \1802 , \1799 , \1801 );
mbuf \mul_17_13/Z[10] ( \1803_Z[10] , \1802 );
mand \U$1/U$149 ( \1804 , \1803_Z[10] , \867 );
mbuf \mul_16_12/A[10] ( \1805_A[10] , \a[10] );
mand \mul_16_12/U$1398 ( \1806 , \1805_A[10] , \892_B[0] );
mand \mul_16_12/U$1383 ( \1807 , \1659_A[9] , \929_B[1] );
mxor \mul_16_12/U$1334 ( \1808 , \1806 , \1807 );
mand \mul_16_12/U$1338 ( \1809 , \1660 , \1661 );
mand \mul_16_12/U$1337 ( \1810 , \1662 , \1665 );
mor \mul_16_12/U$1335 ( \1811 , \1809 , \1810 );
mxor \mul_16_12/U$1331 ( \1812 , \1808 , \1811 );
mand \mul_16_12/U$1294 ( \1813 , \1525_A[8] , \979_B[2] );
mxor \mul_16_12/U$1249 ( \1814 , \1812 , \1813 );
mand \mul_16_12/U$1253 ( \1815 , \1666 , \1667 );
mand \mul_16_12/U$1252 ( \1816 , \1668 , \1671 );
mor \mul_16_12/U$1250 ( \1817 , \1815 , \1816 );
mxor \mul_16_12/U$1246 ( \1818 , \1814 , \1817 );
mand \mul_16_12/U$1202 ( \1819 , \1403_A[7] , \1047_B[3] );
mxor \mul_16_12/U$1161 ( \1820 , \1818 , \1819 );
mand \mul_16_12/U$1165 ( \1821 , \1672 , \1673 );
mand \mul_16_12/U$1164 ( \1822 , \1674 , \1677 );
mor \mul_16_12/U$1162 ( \1823 , \1821 , \1822 );
mxor \mul_16_12/U$1158 ( \1824 , \1820 , \1823 );
mand \mul_16_12/U$1110 ( \1825 , \1293_A[6] , \1127_B[4] );
mxor \mul_16_12/U$1073 ( \1826 , \1824 , \1825 );
mand \mul_16_12/U$1077 ( \1827 , \1678 , \1679 );
mand \mul_16_12/U$1076 ( \1828 , \1680 , \1683 );
mor \mul_16_12/U$1074 ( \1829 , \1827 , \1828 );
mxor \mul_16_12/U$1070 ( \1830 , \1826 , \1829 );
mand \mul_16_12/U$1018 ( \1831 , \1195_A[5] , \1219_B[5] );
mxor \mul_16_12/U$985 ( \1832 , \1830 , \1831 );
mand \mul_16_12/U$989 ( \1833 , \1684 , \1685 );
mand \mul_16_12/U$988 ( \1834 , \1686 , \1689 );
mor \mul_16_12/U$986 ( \1835 , \1833 , \1834 );
mxor \mul_16_12/U$982 ( \1836 , \1832 , \1835 );
mand \mul_16_12/U$926 ( \1837 , \1109_A[4] , \1323_B[6] );
mxor \mul_16_12/U$897 ( \1838 , \1836 , \1837 );
mand \mul_16_12/U$901 ( \1839 , \1690 , \1691 );
mand \mul_16_12/U$900 ( \1840 , \1692 , \1695 );
mor \mul_16_12/U$898 ( \1841 , \1839 , \1840 );
mxor \mul_16_12/U$894 ( \1842 , \1838 , \1841 );
mand \mul_16_12/U$834 ( \1843 , \1035_A[3] , \1439_B[7] );
mxor \mul_16_12/U$809 ( \1844 , \1842 , \1843 );
mand \mul_16_12/U$813 ( \1845 , \1696 , \1697 );
mand \mul_16_12/U$812 ( \1846 , \1698 , \1701 );
mor \mul_16_12/U$810 ( \1847 , \1845 , \1846 );
mxor \mul_16_12/U$806 ( \1848 , \1844 , \1847 );
mand \mul_16_12/U$742 ( \1849 , \973_A[2] , \1567_B[8] );
mxor \mul_16_12/U$721 ( \1850 , \1848 , \1849 );
mand \mul_16_12/U$725 ( \1851 , \1702 , \1703 );
mand \mul_16_12/U$724 ( \1852 , \1704 , \1705 );
mor \mul_16_12/U$722 ( \1853 , \1851 , \1852 );
mxor \mul_16_12/U$718 ( \1854 , \1850 , \1853 );
mand \mul_16_12/U$650 ( \1855 , \927_A[1] , \1707_B[9] );
mxor \mul_16_12/U$633 ( \1856 , \1854 , \1855 );
mand \mul_16_12/U$634 ( \1857 , \1706 , \1708 );
mxor \mul_16_12/U$630 ( \1858 , \1856 , \1857 );
mbuf \mul_16_12/B[10] ( \1859_B[10] , \d[10] );
mand \mul_16_12/U$558 ( \1860 , \891_A[0] , \1859_B[10] );
mxor \mul_16_12/U$542 ( \1861 , \1858 , \1860 );
mbuf \mul_16_12/Z[10] ( \1862_Z[10] , \1861 );
mand \U$1/U$148 ( \1863 , \1862_Z[10] , \865 );
mbuf \add_15_12/A[10] ( \1864_A[10] , \b[10] );
mbuf \add_15_12/B[10] ( \1865_B[10] , \d[10] );
mxor \add_15_12/U$32 ( \1866 , \1864_A[10] , \1865_B[10] );
mand \add_15_12/U$36 ( \1867 , \1712_A[9] , \1713_B[9] );
mand \add_15_12/U$35 ( \1868 , \1713_B[9] , \1718 );
mand \add_15_12/U$34 ( \1869 , \1712_A[9] , \1718 );
mor \add_15_12/U$33 ( \1870 , \1867 , \1868 , \1869 );
mxor \add_15_12/U$31 ( \1871 , \1866 , \1870 );
mbuf \add_15_12/SUM[10] ( \1872_SUM[10] , \1871 );
mand \U$1/U$147 ( \1873 , \1872_SUM[10] , \863 );
mbuf \add_14_12/A[10] ( \1874_A[10] , \a[10] );
mbuf \add_14_12/B[10] ( \1875_B[10] , \c[10] );
mxor \add_14_12/U$32 ( \1876 , \1874_A[10] , \1875_B[10] );
mand \add_14_12/U$36 ( \1877 , \1722_A[9] , \1723_B[9] );
mand \add_14_12/U$35 ( \1878 , \1723_B[9] , \1728 );
mand \add_14_12/U$34 ( \1879 , \1722_A[9] , \1728 );
mor \add_14_12/U$33 ( \1880 , \1877 , \1878 , \1879 );
mxor \add_14_12/U$31 ( \1881 , \1876 , \1880 );
mbuf \add_14_12/SUM[10] ( \1882_SUM[10] , \1881 );
mand \U$1/U$146 ( \1883 , \1882_SUM[10] , \861 );
mand \U$1/U$145 ( \1884 , \d[10] , \859 );
mand \U$1/U$144 ( \1885 , \c[10] , \857 );
mand \U$1/U$143 ( \1886 , \b[10] , \855 );
mand \U$1/U$142 ( \1887 , \a[10] , \853 );
mor \U$1/U$141 ( \1888 , \1737 , \1739 , \1741 , \1743 , \1745 , \1804 , \1863 , \1873 , \1883 , \1884 , \1885 , \1886 , \1887 );
m_DC \n22[11]_g1 ( \1889 , 1'b0 , \876 );
mor \U$5/U$12 ( \1890 , \a[11] , \d[11] );
mand \U$1/U$167 ( \1891 , \1890 , \875 );
mand \U$4/U$12 ( \1892 , \b[11] , \c[11] );
mand \U$1/U$166 ( \1893 , \1892 , \873 );
mor \U$3/U$12 ( \1894 , \a[11] , \b[11] );
mand \U$1/U$165 ( \1895 , \1894 , \871 );
mxor \U$2/U$12 ( \1896 , \c[11] , \d[11] );
mand \U$1/U$164 ( \1897 , \1896 , \869 );
mbuf \mul_17_13/A[11] ( \1898_A[11] , \b[11] );
mand \mul_17_13/U$1397 ( \1899 , \1898_A[11] , \887_B[0] );
mand \mul_17_13/U$1382 ( \1900 , \1746_A[10] , \922_B[1] );
mxor \mul_17_13/U$1329 ( \1901 , \1899 , \1900 );
mand \mul_17_13/U$1333 ( \1902 , \1747 , \1748 );
mand \mul_17_13/U$1332 ( \1903 , \1749 , \1752 );
mor \mul_17_13/U$1330 ( \1904 , \1902 , \1903 );
mxor \mul_17_13/U$1326 ( \1905 , \1901 , \1904 );
mand \mul_17_13/U$1293 ( \1906 , \1606_A[9] , \968_B[2] );
mxor \mul_17_13/U$1244 ( \1907 , \1905 , \1906 );
mand \mul_17_13/U$1248 ( \1908 , \1753 , \1754 );
mand \mul_17_13/U$1247 ( \1909 , \1755 , \1758 );
mor \mul_17_13/U$1245 ( \1910 , \1908 , \1909 );
mxor \mul_17_13/U$1241 ( \1911 , \1907 , \1910 );
mand \mul_17_13/U$1201 ( \1912 , \1478_A[8] , \1030_B[3] );
mxor \mul_17_13/U$1156 ( \1913 , \1911 , \1912 );
mand \mul_17_13/U$1160 ( \1914 , \1759 , \1760 );
mand \mul_17_13/U$1159 ( \1915 , \1761 , \1764 );
mor \mul_17_13/U$1157 ( \1916 , \1914 , \1915 );
mxor \mul_17_13/U$1153 ( \1917 , \1913 , \1916 );
mand \mul_17_13/U$1109 ( \1918 , \1362_A[7] , \1104_B[4] );
mxor \mul_17_13/U$1068 ( \1919 , \1917 , \1918 );
mand \mul_17_13/U$1072 ( \1920 , \1765 , \1766 );
mand \mul_17_13/U$1071 ( \1921 , \1767 , \1770 );
mor \mul_17_13/U$1069 ( \1922 , \1920 , \1921 );
mxor \mul_17_13/U$1065 ( \1923 , \1919 , \1922 );
mand \mul_17_13/U$1017 ( \1924 , \1258_A[6] , \1190_B[5] );
mxor \mul_17_13/U$980 ( \1925 , \1923 , \1924 );
mand \mul_17_13/U$984 ( \1926 , \1771 , \1772 );
mand \mul_17_13/U$983 ( \1927 , \1773 , \1776 );
mor \mul_17_13/U$981 ( \1928 , \1926 , \1927 );
mxor \mul_17_13/U$977 ( \1929 , \1925 , \1928 );
mand \mul_17_13/U$925 ( \1930 , \1166_A[5] , \1288_B[6] );
mxor \mul_17_13/U$892 ( \1931 , \1929 , \1930 );
mand \mul_17_13/U$896 ( \1932 , \1777 , \1778 );
mand \mul_17_13/U$895 ( \1933 , \1779 , \1782 );
mor \mul_17_13/U$893 ( \1934 , \1932 , \1933 );
mxor \mul_17_13/U$889 ( \1935 , \1931 , \1934 );
mand \mul_17_13/U$833 ( \1936 , \1086_A[4] , \1398_B[7] );
mxor \mul_17_13/U$804 ( \1937 , \1935 , \1936 );
mand \mul_17_13/U$808 ( \1938 , \1783 , \1784 );
mand \mul_17_13/U$807 ( \1939 , \1785 , \1788 );
mor \mul_17_13/U$805 ( \1940 , \1938 , \1939 );
mxor \mul_17_13/U$801 ( \1941 , \1937 , \1940 );
mand \mul_17_13/U$741 ( \1942 , \1018_A[3] , \1520_B[8] );
mxor \mul_17_13/U$716 ( \1943 , \1941 , \1942 );
mand \mul_17_13/U$720 ( \1944 , \1789 , \1790 );
mand \mul_17_13/U$719 ( \1945 , \1791 , \1794 );
mor \mul_17_13/U$717 ( \1946 , \1944 , \1945 );
mxor \mul_17_13/U$713 ( \1947 , \1943 , \1946 );
mand \mul_17_13/U$649 ( \1948 , \962_A[2] , \1654_B[9] );
mxor \mul_17_13/U$628 ( \1949 , \1947 , \1948 );
mand \mul_17_13/U$632 ( \1950 , \1795 , \1796 );
mand \mul_17_13/U$631 ( \1951 , \1797 , \1798 );
mor \mul_17_13/U$629 ( \1952 , \1950 , \1951 );
mxor \mul_17_13/U$625 ( \1953 , \1949 , \1952 );
mand \mul_17_13/U$557 ( \1954 , \920_A[1] , \1800_B[10] );
mxor \mul_17_13/U$540 ( \1955 , \1953 , \1954 );
mand \mul_17_13/U$541 ( \1956 , \1799 , \1801 );
mxor \mul_17_13/U$537 ( \1957 , \1955 , \1956 );
mbuf \mul_17_13/B[11] ( \1958_B[11] , \c[11] );
mand \mul_17_13/U$465 ( \1959 , \886_A[0] , \1958_B[11] );
mxor \mul_17_13/U$449 ( \1960 , \1957 , \1959 );
mbuf \mul_17_13/Z[11] ( \1961_Z[11] , \1960 );
mand \U$1/U$163 ( \1962 , \1961_Z[11] , \867 );
mbuf \mul_16_12/A[11] ( \1963_A[11] , \a[11] );
mand \mul_16_12/U$1397 ( \1964 , \1963_A[11] , \892_B[0] );
mand \mul_16_12/U$1382 ( \1965 , \1805_A[10] , \929_B[1] );
mxor \mul_16_12/U$1329 ( \1966 , \1964 , \1965 );
mand \mul_16_12/U$1333 ( \1967 , \1806 , \1807 );
mand \mul_16_12/U$1332 ( \1968 , \1808 , \1811 );
mor \mul_16_12/U$1330 ( \1969 , \1967 , \1968 );
mxor \mul_16_12/U$1326 ( \1970 , \1966 , \1969 );
mand \mul_16_12/U$1293 ( \1971 , \1659_A[9] , \979_B[2] );
mxor \mul_16_12/U$1244 ( \1972 , \1970 , \1971 );
mand \mul_16_12/U$1248 ( \1973 , \1812 , \1813 );
mand \mul_16_12/U$1247 ( \1974 , \1814 , \1817 );
mor \mul_16_12/U$1245 ( \1975 , \1973 , \1974 );
mxor \mul_16_12/U$1241 ( \1976 , \1972 , \1975 );
mand \mul_16_12/U$1201 ( \1977 , \1525_A[8] , \1047_B[3] );
mxor \mul_16_12/U$1156 ( \1978 , \1976 , \1977 );
mand \mul_16_12/U$1160 ( \1979 , \1818 , \1819 );
mand \mul_16_12/U$1159 ( \1980 , \1820 , \1823 );
mor \mul_16_12/U$1157 ( \1981 , \1979 , \1980 );
mxor \mul_16_12/U$1153 ( \1982 , \1978 , \1981 );
mand \mul_16_12/U$1109 ( \1983 , \1403_A[7] , \1127_B[4] );
mxor \mul_16_12/U$1068 ( \1984 , \1982 , \1983 );
mand \mul_16_12/U$1072 ( \1985 , \1824 , \1825 );
mand \mul_16_12/U$1071 ( \1986 , \1826 , \1829 );
mor \mul_16_12/U$1069 ( \1987 , \1985 , \1986 );
mxor \mul_16_12/U$1065 ( \1988 , \1984 , \1987 );
mand \mul_16_12/U$1017 ( \1989 , \1293_A[6] , \1219_B[5] );
mxor \mul_16_12/U$980 ( \1990 , \1988 , \1989 );
mand \mul_16_12/U$984 ( \1991 , \1830 , \1831 );
mand \mul_16_12/U$983 ( \1992 , \1832 , \1835 );
mor \mul_16_12/U$981 ( \1993 , \1991 , \1992 );
mxor \mul_16_12/U$977 ( \1994 , \1990 , \1993 );
mand \mul_16_12/U$925 ( \1995 , \1195_A[5] , \1323_B[6] );
mxor \mul_16_12/U$892 ( \1996 , \1994 , \1995 );
mand \mul_16_12/U$896 ( \1997 , \1836 , \1837 );
mand \mul_16_12/U$895 ( \1998 , \1838 , \1841 );
mor \mul_16_12/U$893 ( \1999 , \1997 , \1998 );
mxor \mul_16_12/U$889 ( \2000 , \1996 , \1999 );
mand \mul_16_12/U$833 ( \2001 , \1109_A[4] , \1439_B[7] );
mxor \mul_16_12/U$804 ( \2002 , \2000 , \2001 );
mand \mul_16_12/U$808 ( \2003 , \1842 , \1843 );
mand \mul_16_12/U$807 ( \2004 , \1844 , \1847 );
mor \mul_16_12/U$805 ( \2005 , \2003 , \2004 );
mxor \mul_16_12/U$801 ( \2006 , \2002 , \2005 );
mand \mul_16_12/U$741 ( \2007 , \1035_A[3] , \1567_B[8] );
mxor \mul_16_12/U$716 ( \2008 , \2006 , \2007 );
mand \mul_16_12/U$720 ( \2009 , \1848 , \1849 );
mand \mul_16_12/U$719 ( \2010 , \1850 , \1853 );
mor \mul_16_12/U$717 ( \2011 , \2009 , \2010 );
mxor \mul_16_12/U$713 ( \2012 , \2008 , \2011 );
mand \mul_16_12/U$649 ( \2013 , \973_A[2] , \1707_B[9] );
mxor \mul_16_12/U$628 ( \2014 , \2012 , \2013 );
mand \mul_16_12/U$632 ( \2015 , \1854 , \1855 );
mand \mul_16_12/U$631 ( \2016 , \1856 , \1857 );
mor \mul_16_12/U$629 ( \2017 , \2015 , \2016 );
mxor \mul_16_12/U$625 ( \2018 , \2014 , \2017 );
mand \mul_16_12/U$557 ( \2019 , \927_A[1] , \1859_B[10] );
mxor \mul_16_12/U$540 ( \2020 , \2018 , \2019 );
mand \mul_16_12/U$541 ( \2021 , \1858 , \1860 );
mxor \mul_16_12/U$537 ( \2022 , \2020 , \2021 );
mbuf \mul_16_12/B[11] ( \2023_B[11] , \d[11] );
mand \mul_16_12/U$465 ( \2024 , \891_A[0] , \2023_B[11] );
mxor \mul_16_12/U$449 ( \2025 , \2022 , \2024 );
mbuf \mul_16_12/Z[11] ( \2026_Z[11] , \2025 );
mand \U$1/U$162 ( \2027 , \2026_Z[11] , \865 );
mbuf \add_15_12/A[11] ( \2028_A[11] , \b[11] );
mbuf \add_15_12/B[11] ( \2029_B[11] , \d[11] );
mxor \add_15_12/U$26 ( \2030 , \2028_A[11] , \2029_B[11] );
mand \add_15_12/U$30 ( \2031 , \1864_A[10] , \1865_B[10] );
mand \add_15_12/U$29 ( \2032 , \1865_B[10] , \1870 );
mand \add_15_12/U$28 ( \2033 , \1864_A[10] , \1870 );
mor \add_15_12/U$27 ( \2034 , \2031 , \2032 , \2033 );
mxor \add_15_12/U$25 ( \2035 , \2030 , \2034 );
mbuf \add_15_12/SUM[11] ( \2036_SUM[11] , \2035 );
mand \U$1/U$161 ( \2037 , \2036_SUM[11] , \863 );
mbuf \add_14_12/A[11] ( \2038_A[11] , \a[11] );
mbuf \add_14_12/B[11] ( \2039_B[11] , \c[11] );
mxor \add_14_12/U$26 ( \2040 , \2038_A[11] , \2039_B[11] );
mand \add_14_12/U$30 ( \2041 , \1874_A[10] , \1875_B[10] );
mand \add_14_12/U$29 ( \2042 , \1875_B[10] , \1880 );
mand \add_14_12/U$28 ( \2043 , \1874_A[10] , \1880 );
mor \add_14_12/U$27 ( \2044 , \2041 , \2042 , \2043 );
mxor \add_14_12/U$25 ( \2045 , \2040 , \2044 );
mbuf \add_14_12/SUM[11] ( \2046_SUM[11] , \2045 );
mand \U$1/U$160 ( \2047 , \2046_SUM[11] , \861 );
mand \U$1/U$159 ( \2048 , \d[11] , \859 );
mand \U$1/U$158 ( \2049 , \c[11] , \857 );
mand \U$1/U$157 ( \2050 , \b[11] , \855 );
mand \U$1/U$156 ( \2051 , \a[11] , \853 );
mor \U$1/U$155 ( \2052 , \1889 , \1891 , \1893 , \1895 , \1897 , \1962 , \2027 , \2037 , \2047 , \2048 , \2049 , \2050 , \2051 );
m_DC \n22[12]_g1 ( \2053 , 1'b0 , \876 );
mor \U$5/U$13 ( \2054 , \a[12] , \d[12] );
mand \U$1/U$181 ( \2055 , \2054 , \875 );
mand \U$4/U$13 ( \2056 , \b[12] , \c[12] );
mand \U$1/U$180 ( \2057 , \2056 , \873 );
mor \U$3/U$13 ( \2058 , \a[12] , \b[12] );
mand \U$1/U$179 ( \2059 , \2058 , \871 );
mxor \U$2/U$13 ( \2060 , \c[12] , \d[12] );
mand \U$1/U$178 ( \2061 , \2060 , \869 );
mbuf \mul_17_13/A[12] ( \2062_A[12] , \b[12] );
mand \mul_17_13/U$1396 ( \2063 , \2062_A[12] , \887_B[0] );
mand \mul_17_13/U$1381 ( \2064 , \1898_A[11] , \922_B[1] );
mxor \mul_17_13/U$1324 ( \2065 , \2063 , \2064 );
mand \mul_17_13/U$1328 ( \2066 , \1899 , \1900 );
mand \mul_17_13/U$1327 ( \2067 , \1901 , \1904 );
mor \mul_17_13/U$1325 ( \2068 , \2066 , \2067 );
mxor \mul_17_13/U$1321 ( \2069 , \2065 , \2068 );
mand \mul_17_13/U$1292 ( \2070 , \1746_A[10] , \968_B[2] );
mxor \mul_17_13/U$1239 ( \2071 , \2069 , \2070 );
mand \mul_17_13/U$1243 ( \2072 , \1905 , \1906 );
mand \mul_17_13/U$1242 ( \2073 , \1907 , \1910 );
mor \mul_17_13/U$1240 ( \2074 , \2072 , \2073 );
mxor \mul_17_13/U$1236 ( \2075 , \2071 , \2074 );
mand \mul_17_13/U$1200 ( \2076 , \1606_A[9] , \1030_B[3] );
mxor \mul_17_13/U$1151 ( \2077 , \2075 , \2076 );
mand \mul_17_13/U$1155 ( \2078 , \1911 , \1912 );
mand \mul_17_13/U$1154 ( \2079 , \1913 , \1916 );
mor \mul_17_13/U$1152 ( \2080 , \2078 , \2079 );
mxor \mul_17_13/U$1148 ( \2081 , \2077 , \2080 );
mand \mul_17_13/U$1108 ( \2082 , \1478_A[8] , \1104_B[4] );
mxor \mul_17_13/U$1063 ( \2083 , \2081 , \2082 );
mand \mul_17_13/U$1067 ( \2084 , \1917 , \1918 );
mand \mul_17_13/U$1066 ( \2085 , \1919 , \1922 );
mor \mul_17_13/U$1064 ( \2086 , \2084 , \2085 );
mxor \mul_17_13/U$1060 ( \2087 , \2083 , \2086 );
mand \mul_17_13/U$1016 ( \2088 , \1362_A[7] , \1190_B[5] );
mxor \mul_17_13/U$975 ( \2089 , \2087 , \2088 );
mand \mul_17_13/U$979 ( \2090 , \1923 , \1924 );
mand \mul_17_13/U$978 ( \2091 , \1925 , \1928 );
mor \mul_17_13/U$976 ( \2092 , \2090 , \2091 );
mxor \mul_17_13/U$972 ( \2093 , \2089 , \2092 );
mand \mul_17_13/U$924 ( \2094 , \1258_A[6] , \1288_B[6] );
mxor \mul_17_13/U$887 ( \2095 , \2093 , \2094 );
mand \mul_17_13/U$891 ( \2096 , \1929 , \1930 );
mand \mul_17_13/U$890 ( \2097 , \1931 , \1934 );
mor \mul_17_13/U$888 ( \2098 , \2096 , \2097 );
mxor \mul_17_13/U$884 ( \2099 , \2095 , \2098 );
mand \mul_17_13/U$832 ( \2100 , \1166_A[5] , \1398_B[7] );
mxor \mul_17_13/U$799 ( \2101 , \2099 , \2100 );
mand \mul_17_13/U$803 ( \2102 , \1935 , \1936 );
mand \mul_17_13/U$802 ( \2103 , \1937 , \1940 );
mor \mul_17_13/U$800 ( \2104 , \2102 , \2103 );
mxor \mul_17_13/U$796 ( \2105 , \2101 , \2104 );
mand \mul_17_13/U$740 ( \2106 , \1086_A[4] , \1520_B[8] );
mxor \mul_17_13/U$711 ( \2107 , \2105 , \2106 );
mand \mul_17_13/U$715 ( \2108 , \1941 , \1942 );
mand \mul_17_13/U$714 ( \2109 , \1943 , \1946 );
mor \mul_17_13/U$712 ( \2110 , \2108 , \2109 );
mxor \mul_17_13/U$708 ( \2111 , \2107 , \2110 );
mand \mul_17_13/U$648 ( \2112 , \1018_A[3] , \1654_B[9] );
mxor \mul_17_13/U$623 ( \2113 , \2111 , \2112 );
mand \mul_17_13/U$627 ( \2114 , \1947 , \1948 );
mand \mul_17_13/U$626 ( \2115 , \1949 , \1952 );
mor \mul_17_13/U$624 ( \2116 , \2114 , \2115 );
mxor \mul_17_13/U$620 ( \2117 , \2113 , \2116 );
mand \mul_17_13/U$556 ( \2118 , \962_A[2] , \1800_B[10] );
mxor \mul_17_13/U$535 ( \2119 , \2117 , \2118 );
mand \mul_17_13/U$539 ( \2120 , \1953 , \1954 );
mand \mul_17_13/U$538 ( \2121 , \1955 , \1956 );
mor \mul_17_13/U$536 ( \2122 , \2120 , \2121 );
mxor \mul_17_13/U$532 ( \2123 , \2119 , \2122 );
mand \mul_17_13/U$464 ( \2124 , \920_A[1] , \1958_B[11] );
mxor \mul_17_13/U$447 ( \2125 , \2123 , \2124 );
mand \mul_17_13/U$448 ( \2126 , \1957 , \1959 );
mxor \mul_17_13/U$444 ( \2127 , \2125 , \2126 );
mbuf \mul_17_13/B[12] ( \2128_B[12] , \c[12] );
mand \mul_17_13/U$372 ( \2129 , \886_A[0] , \2128_B[12] );
mxor \mul_17_13/U$356 ( \2130 , \2127 , \2129 );
mbuf \mul_17_13/Z[12] ( \2131_Z[12] , \2130 );
mand \U$1/U$177 ( \2132 , \2131_Z[12] , \867 );
mbuf \mul_16_12/A[12] ( \2133_A[12] , \a[12] );
mand \mul_16_12/U$1396 ( \2134 , \2133_A[12] , \892_B[0] );
mand \mul_16_12/U$1381 ( \2135 , \1963_A[11] , \929_B[1] );
mxor \mul_16_12/U$1324 ( \2136 , \2134 , \2135 );
mand \mul_16_12/U$1328 ( \2137 , \1964 , \1965 );
mand \mul_16_12/U$1327 ( \2138 , \1966 , \1969 );
mor \mul_16_12/U$1325 ( \2139 , \2137 , \2138 );
mxor \mul_16_12/U$1321 ( \2140 , \2136 , \2139 );
mand \mul_16_12/U$1292 ( \2141 , \1805_A[10] , \979_B[2] );
mxor \mul_16_12/U$1239 ( \2142 , \2140 , \2141 );
mand \mul_16_12/U$1243 ( \2143 , \1970 , \1971 );
mand \mul_16_12/U$1242 ( \2144 , \1972 , \1975 );
mor \mul_16_12/U$1240 ( \2145 , \2143 , \2144 );
mxor \mul_16_12/U$1236 ( \2146 , \2142 , \2145 );
mand \mul_16_12/U$1200 ( \2147 , \1659_A[9] , \1047_B[3] );
mxor \mul_16_12/U$1151 ( \2148 , \2146 , \2147 );
mand \mul_16_12/U$1155 ( \2149 , \1976 , \1977 );
mand \mul_16_12/U$1154 ( \2150 , \1978 , \1981 );
mor \mul_16_12/U$1152 ( \2151 , \2149 , \2150 );
mxor \mul_16_12/U$1148 ( \2152 , \2148 , \2151 );
mand \mul_16_12/U$1108 ( \2153 , \1525_A[8] , \1127_B[4] );
mxor \mul_16_12/U$1063 ( \2154 , \2152 , \2153 );
mand \mul_16_12/U$1067 ( \2155 , \1982 , \1983 );
mand \mul_16_12/U$1066 ( \2156 , \1984 , \1987 );
mor \mul_16_12/U$1064 ( \2157 , \2155 , \2156 );
mxor \mul_16_12/U$1060 ( \2158 , \2154 , \2157 );
mand \mul_16_12/U$1016 ( \2159 , \1403_A[7] , \1219_B[5] );
mxor \mul_16_12/U$975 ( \2160 , \2158 , \2159 );
mand \mul_16_12/U$979 ( \2161 , \1988 , \1989 );
mand \mul_16_12/U$978 ( \2162 , \1990 , \1993 );
mor \mul_16_12/U$976 ( \2163 , \2161 , \2162 );
mxor \mul_16_12/U$972 ( \2164 , \2160 , \2163 );
mand \mul_16_12/U$924 ( \2165 , \1293_A[6] , \1323_B[6] );
mxor \mul_16_12/U$887 ( \2166 , \2164 , \2165 );
mand \mul_16_12/U$891 ( \2167 , \1994 , \1995 );
mand \mul_16_12/U$890 ( \2168 , \1996 , \1999 );
mor \mul_16_12/U$888 ( \2169 , \2167 , \2168 );
mxor \mul_16_12/U$884 ( \2170 , \2166 , \2169 );
mand \mul_16_12/U$832 ( \2171 , \1195_A[5] , \1439_B[7] );
mxor \mul_16_12/U$799 ( \2172 , \2170 , \2171 );
mand \mul_16_12/U$803 ( \2173 , \2000 , \2001 );
mand \mul_16_12/U$802 ( \2174 , \2002 , \2005 );
mor \mul_16_12/U$800 ( \2175 , \2173 , \2174 );
mxor \mul_16_12/U$796 ( \2176 , \2172 , \2175 );
mand \mul_16_12/U$740 ( \2177 , \1109_A[4] , \1567_B[8] );
mxor \mul_16_12/U$711 ( \2178 , \2176 , \2177 );
mand \mul_16_12/U$715 ( \2179 , \2006 , \2007 );
mand \mul_16_12/U$714 ( \2180 , \2008 , \2011 );
mor \mul_16_12/U$712 ( \2181 , \2179 , \2180 );
mxor \mul_16_12/U$708 ( \2182 , \2178 , \2181 );
mand \mul_16_12/U$648 ( \2183 , \1035_A[3] , \1707_B[9] );
mxor \mul_16_12/U$623 ( \2184 , \2182 , \2183 );
mand \mul_16_12/U$627 ( \2185 , \2012 , \2013 );
mand \mul_16_12/U$626 ( \2186 , \2014 , \2017 );
mor \mul_16_12/U$624 ( \2187 , \2185 , \2186 );
mxor \mul_16_12/U$620 ( \2188 , \2184 , \2187 );
mand \mul_16_12/U$556 ( \2189 , \973_A[2] , \1859_B[10] );
mxor \mul_16_12/U$535 ( \2190 , \2188 , \2189 );
mand \mul_16_12/U$539 ( \2191 , \2018 , \2019 );
mand \mul_16_12/U$538 ( \2192 , \2020 , \2021 );
mor \mul_16_12/U$536 ( \2193 , \2191 , \2192 );
mxor \mul_16_12/U$532 ( \2194 , \2190 , \2193 );
mand \mul_16_12/U$464 ( \2195 , \927_A[1] , \2023_B[11] );
mxor \mul_16_12/U$447 ( \2196 , \2194 , \2195 );
mand \mul_16_12/U$448 ( \2197 , \2022 , \2024 );
mxor \mul_16_12/U$444 ( \2198 , \2196 , \2197 );
mbuf \mul_16_12/B[12] ( \2199_B[12] , \d[12] );
mand \mul_16_12/U$372 ( \2200 , \891_A[0] , \2199_B[12] );
mxor \mul_16_12/U$356 ( \2201 , \2198 , \2200 );
mbuf \mul_16_12/Z[12] ( \2202_Z[12] , \2201 );
mand \U$1/U$176 ( \2203 , \2202_Z[12] , \865 );
mbuf \add_15_12/A[12] ( \2204_A[12] , \b[12] );
mbuf \add_15_12/B[12] ( \2205_B[12] , \d[12] );
mxor \add_15_12/U$20 ( \2206 , \2204_A[12] , \2205_B[12] );
mand \add_15_12/U$24 ( \2207 , \2028_A[11] , \2029_B[11] );
mand \add_15_12/U$23 ( \2208 , \2029_B[11] , \2034 );
mand \add_15_12/U$22 ( \2209 , \2028_A[11] , \2034 );
mor \add_15_12/U$21 ( \2210 , \2207 , \2208 , \2209 );
mxor \add_15_12/U$19 ( \2211 , \2206 , \2210 );
mbuf \add_15_12/SUM[12] ( \2212_SUM[12] , \2211 );
mand \U$1/U$175 ( \2213 , \2212_SUM[12] , \863 );
mbuf \add_14_12/A[12] ( \2214_A[12] , \a[12] );
mbuf \add_14_12/B[12] ( \2215_B[12] , \c[12] );
mxor \add_14_12/U$20 ( \2216 , \2214_A[12] , \2215_B[12] );
mand \add_14_12/U$24 ( \2217 , \2038_A[11] , \2039_B[11] );
mand \add_14_12/U$23 ( \2218 , \2039_B[11] , \2044 );
mand \add_14_12/U$22 ( \2219 , \2038_A[11] , \2044 );
mor \add_14_12/U$21 ( \2220 , \2217 , \2218 , \2219 );
mxor \add_14_12/U$19 ( \2221 , \2216 , \2220 );
mbuf \add_14_12/SUM[12] ( \2222_SUM[12] , \2221 );
mand \U$1/U$174 ( \2223 , \2222_SUM[12] , \861 );
mand \U$1/U$173 ( \2224 , \d[12] , \859 );
mand \U$1/U$172 ( \2225 , \c[12] , \857 );
mand \U$1/U$171 ( \2226 , \b[12] , \855 );
mand \U$1/U$170 ( \2227 , \a[12] , \853 );
mor \U$1/U$169 ( \2228 , \2053 , \2055 , \2057 , \2059 , \2061 , \2132 , \2203 , \2213 , \2223 , \2224 , \2225 , \2226 , \2227 );
m_DC \n22[13]_g1 ( \2229 , 1'b0 , \876 );
mor \U$5/U$14 ( \2230 , \a[13] , \d[13] );
mand \U$1/U$195 ( \2231 , \2230 , \875 );
mand \U$4/U$14 ( \2232 , \b[13] , \c[13] );
mand \U$1/U$194 ( \2233 , \2232 , \873 );
mor \U$3/U$14 ( \2234 , \a[13] , \b[13] );
mand \U$1/U$193 ( \2235 , \2234 , \871 );
mxor \U$2/U$14 ( \2236 , \c[13] , \d[13] );
mand \U$1/U$192 ( \2237 , \2236 , \869 );
mbuf \mul_17_13/A[13] ( \2238_A[13] , \b[13] );
mand \mul_17_13/U$1395 ( \2239 , \2238_A[13] , \887_B[0] );
mand \mul_17_13/U$1380 ( \2240 , \2062_A[12] , \922_B[1] );
mxor \mul_17_13/U$1319 ( \2241 , \2239 , \2240 );
mand \mul_17_13/U$1323 ( \2242 , \2063 , \2064 );
mand \mul_17_13/U$1322 ( \2243 , \2065 , \2068 );
mor \mul_17_13/U$1320 ( \2244 , \2242 , \2243 );
mxor \mul_17_13/U$1316 ( \2245 , \2241 , \2244 );
mand \mul_17_13/U$1291 ( \2246 , \1898_A[11] , \968_B[2] );
mxor \mul_17_13/U$1234 ( \2247 , \2245 , \2246 );
mand \mul_17_13/U$1238 ( \2248 , \2069 , \2070 );
mand \mul_17_13/U$1237 ( \2249 , \2071 , \2074 );
mor \mul_17_13/U$1235 ( \2250 , \2248 , \2249 );
mxor \mul_17_13/U$1231 ( \2251 , \2247 , \2250 );
mand \mul_17_13/U$1199 ( \2252 , \1746_A[10] , \1030_B[3] );
mxor \mul_17_13/U$1146 ( \2253 , \2251 , \2252 );
mand \mul_17_13/U$1150 ( \2254 , \2075 , \2076 );
mand \mul_17_13/U$1149 ( \2255 , \2077 , \2080 );
mor \mul_17_13/U$1147 ( \2256 , \2254 , \2255 );
mxor \mul_17_13/U$1143 ( \2257 , \2253 , \2256 );
mand \mul_17_13/U$1107 ( \2258 , \1606_A[9] , \1104_B[4] );
mxor \mul_17_13/U$1058 ( \2259 , \2257 , \2258 );
mand \mul_17_13/U$1062 ( \2260 , \2081 , \2082 );
mand \mul_17_13/U$1061 ( \2261 , \2083 , \2086 );
mor \mul_17_13/U$1059 ( \2262 , \2260 , \2261 );
mxor \mul_17_13/U$1055 ( \2263 , \2259 , \2262 );
mand \mul_17_13/U$1015 ( \2264 , \1478_A[8] , \1190_B[5] );
mxor \mul_17_13/U$970 ( \2265 , \2263 , \2264 );
mand \mul_17_13/U$974 ( \2266 , \2087 , \2088 );
mand \mul_17_13/U$973 ( \2267 , \2089 , \2092 );
mor \mul_17_13/U$971 ( \2268 , \2266 , \2267 );
mxor \mul_17_13/U$967 ( \2269 , \2265 , \2268 );
mand \mul_17_13/U$923 ( \2270 , \1362_A[7] , \1288_B[6] );
mxor \mul_17_13/U$882 ( \2271 , \2269 , \2270 );
mand \mul_17_13/U$886 ( \2272 , \2093 , \2094 );
mand \mul_17_13/U$885 ( \2273 , \2095 , \2098 );
mor \mul_17_13/U$883 ( \2274 , \2272 , \2273 );
mxor \mul_17_13/U$879 ( \2275 , \2271 , \2274 );
mand \mul_17_13/U$831 ( \2276 , \1258_A[6] , \1398_B[7] );
mxor \mul_17_13/U$794 ( \2277 , \2275 , \2276 );
mand \mul_17_13/U$798 ( \2278 , \2099 , \2100 );
mand \mul_17_13/U$797 ( \2279 , \2101 , \2104 );
mor \mul_17_13/U$795 ( \2280 , \2278 , \2279 );
mxor \mul_17_13/U$791 ( \2281 , \2277 , \2280 );
mand \mul_17_13/U$739 ( \2282 , \1166_A[5] , \1520_B[8] );
mxor \mul_17_13/U$706 ( \2283 , \2281 , \2282 );
mand \mul_17_13/U$710 ( \2284 , \2105 , \2106 );
mand \mul_17_13/U$709 ( \2285 , \2107 , \2110 );
mor \mul_17_13/U$707 ( \2286 , \2284 , \2285 );
mxor \mul_17_13/U$703 ( \2287 , \2283 , \2286 );
mand \mul_17_13/U$647 ( \2288 , \1086_A[4] , \1654_B[9] );
mxor \mul_17_13/U$618 ( \2289 , \2287 , \2288 );
mand \mul_17_13/U$622 ( \2290 , \2111 , \2112 );
mand \mul_17_13/U$621 ( \2291 , \2113 , \2116 );
mor \mul_17_13/U$619 ( \2292 , \2290 , \2291 );
mxor \mul_17_13/U$615 ( \2293 , \2289 , \2292 );
mand \mul_17_13/U$555 ( \2294 , \1018_A[3] , \1800_B[10] );
mxor \mul_17_13/U$530 ( \2295 , \2293 , \2294 );
mand \mul_17_13/U$534 ( \2296 , \2117 , \2118 );
mand \mul_17_13/U$533 ( \2297 , \2119 , \2122 );
mor \mul_17_13/U$531 ( \2298 , \2296 , \2297 );
mxor \mul_17_13/U$527 ( \2299 , \2295 , \2298 );
mand \mul_17_13/U$463 ( \2300 , \962_A[2] , \1958_B[11] );
mxor \mul_17_13/U$442 ( \2301 , \2299 , \2300 );
mand \mul_17_13/U$446 ( \2302 , \2123 , \2124 );
mand \mul_17_13/U$445 ( \2303 , \2125 , \2126 );
mor \mul_17_13/U$443 ( \2304 , \2302 , \2303 );
mxor \mul_17_13/U$439 ( \2305 , \2301 , \2304 );
mand \mul_17_13/U$371 ( \2306 , \920_A[1] , \2128_B[12] );
mxor \mul_17_13/U$354 ( \2307 , \2305 , \2306 );
mand \mul_17_13/U$355 ( \2308 , \2127 , \2129 );
mxor \mul_17_13/U$351 ( \2309 , \2307 , \2308 );
mbuf \mul_17_13/B[13] ( \2310_B[13] , \c[13] );
mand \mul_17_13/U$279 ( \2311 , \886_A[0] , \2310_B[13] );
mxor \mul_17_13/U$263 ( \2312 , \2309 , \2311 );
mbuf \mul_17_13/Z[13] ( \2313_Z[13] , \2312 );
mand \U$1/U$191 ( \2314 , \2313_Z[13] , \867 );
mbuf \mul_16_12/A[13] ( \2315_A[13] , \a[13] );
mand \mul_16_12/U$1395 ( \2316 , \2315_A[13] , \892_B[0] );
mand \mul_16_12/U$1380 ( \2317 , \2133_A[12] , \929_B[1] );
mxor \mul_16_12/U$1319 ( \2318 , \2316 , \2317 );
mand \mul_16_12/U$1323 ( \2319 , \2134 , \2135 );
mand \mul_16_12/U$1322 ( \2320 , \2136 , \2139 );
mor \mul_16_12/U$1320 ( \2321 , \2319 , \2320 );
mxor \mul_16_12/U$1316 ( \2322 , \2318 , \2321 );
mand \mul_16_12/U$1291 ( \2323 , \1963_A[11] , \979_B[2] );
mxor \mul_16_12/U$1234 ( \2324 , \2322 , \2323 );
mand \mul_16_12/U$1238 ( \2325 , \2140 , \2141 );
mand \mul_16_12/U$1237 ( \2326 , \2142 , \2145 );
mor \mul_16_12/U$1235 ( \2327 , \2325 , \2326 );
mxor \mul_16_12/U$1231 ( \2328 , \2324 , \2327 );
mand \mul_16_12/U$1199 ( \2329 , \1805_A[10] , \1047_B[3] );
mxor \mul_16_12/U$1146 ( \2330 , \2328 , \2329 );
mand \mul_16_12/U$1150 ( \2331 , \2146 , \2147 );
mand \mul_16_12/U$1149 ( \2332 , \2148 , \2151 );
mor \mul_16_12/U$1147 ( \2333 , \2331 , \2332 );
mxor \mul_16_12/U$1143 ( \2334 , \2330 , \2333 );
mand \mul_16_12/U$1107 ( \2335 , \1659_A[9] , \1127_B[4] );
mxor \mul_16_12/U$1058 ( \2336 , \2334 , \2335 );
mand \mul_16_12/U$1062 ( \2337 , \2152 , \2153 );
mand \mul_16_12/U$1061 ( \2338 , \2154 , \2157 );
mor \mul_16_12/U$1059 ( \2339 , \2337 , \2338 );
mxor \mul_16_12/U$1055 ( \2340 , \2336 , \2339 );
mand \mul_16_12/U$1015 ( \2341 , \1525_A[8] , \1219_B[5] );
mxor \mul_16_12/U$970 ( \2342 , \2340 , \2341 );
mand \mul_16_12/U$974 ( \2343 , \2158 , \2159 );
mand \mul_16_12/U$973 ( \2344 , \2160 , \2163 );
mor \mul_16_12/U$971 ( \2345 , \2343 , \2344 );
mxor \mul_16_12/U$967 ( \2346 , \2342 , \2345 );
mand \mul_16_12/U$923 ( \2347 , \1403_A[7] , \1323_B[6] );
mxor \mul_16_12/U$882 ( \2348 , \2346 , \2347 );
mand \mul_16_12/U$886 ( \2349 , \2164 , \2165 );
mand \mul_16_12/U$885 ( \2350 , \2166 , \2169 );
mor \mul_16_12/U$883 ( \2351 , \2349 , \2350 );
mxor \mul_16_12/U$879 ( \2352 , \2348 , \2351 );
mand \mul_16_12/U$831 ( \2353 , \1293_A[6] , \1439_B[7] );
mxor \mul_16_12/U$794 ( \2354 , \2352 , \2353 );
mand \mul_16_12/U$798 ( \2355 , \2170 , \2171 );
mand \mul_16_12/U$797 ( \2356 , \2172 , \2175 );
mor \mul_16_12/U$795 ( \2357 , \2355 , \2356 );
mxor \mul_16_12/U$791 ( \2358 , \2354 , \2357 );
mand \mul_16_12/U$739 ( \2359 , \1195_A[5] , \1567_B[8] );
mxor \mul_16_12/U$706 ( \2360 , \2358 , \2359 );
mand \mul_16_12/U$710 ( \2361 , \2176 , \2177 );
mand \mul_16_12/U$709 ( \2362 , \2178 , \2181 );
mor \mul_16_12/U$707 ( \2363 , \2361 , \2362 );
mxor \mul_16_12/U$703 ( \2364 , \2360 , \2363 );
mand \mul_16_12/U$647 ( \2365 , \1109_A[4] , \1707_B[9] );
mxor \mul_16_12/U$618 ( \2366 , \2364 , \2365 );
mand \mul_16_12/U$622 ( \2367 , \2182 , \2183 );
mand \mul_16_12/U$621 ( \2368 , \2184 , \2187 );
mor \mul_16_12/U$619 ( \2369 , \2367 , \2368 );
mxor \mul_16_12/U$615 ( \2370 , \2366 , \2369 );
mand \mul_16_12/U$555 ( \2371 , \1035_A[3] , \1859_B[10] );
mxor \mul_16_12/U$530 ( \2372 , \2370 , \2371 );
mand \mul_16_12/U$534 ( \2373 , \2188 , \2189 );
mand \mul_16_12/U$533 ( \2374 , \2190 , \2193 );
mor \mul_16_12/U$531 ( \2375 , \2373 , \2374 );
mxor \mul_16_12/U$527 ( \2376 , \2372 , \2375 );
mand \mul_16_12/U$463 ( \2377 , \973_A[2] , \2023_B[11] );
mxor \mul_16_12/U$442 ( \2378 , \2376 , \2377 );
mand \mul_16_12/U$446 ( \2379 , \2194 , \2195 );
mand \mul_16_12/U$445 ( \2380 , \2196 , \2197 );
mor \mul_16_12/U$443 ( \2381 , \2379 , \2380 );
mxor \mul_16_12/U$439 ( \2382 , \2378 , \2381 );
mand \mul_16_12/U$371 ( \2383 , \927_A[1] , \2199_B[12] );
mxor \mul_16_12/U$354 ( \2384 , \2382 , \2383 );
mand \mul_16_12/U$355 ( \2385 , \2198 , \2200 );
mxor \mul_16_12/U$351 ( \2386 , \2384 , \2385 );
mbuf \mul_16_12/B[13] ( \2387_B[13] , \d[13] );
mand \mul_16_12/U$279 ( \2388 , \891_A[0] , \2387_B[13] );
mxor \mul_16_12/U$263 ( \2389 , \2386 , \2388 );
mbuf \mul_16_12/Z[13] ( \2390_Z[13] , \2389 );
mand \U$1/U$190 ( \2391 , \2390_Z[13] , \865 );
mbuf \add_15_12/A[13] ( \2392_A[13] , \b[13] );
mbuf \add_15_12/B[13] ( \2393_B[13] , \d[13] );
mxor \add_15_12/U$14 ( \2394 , \2392_A[13] , \2393_B[13] );
mand \add_15_12/U$18 ( \2395 , \2204_A[12] , \2205_B[12] );
mand \add_15_12/U$17 ( \2396 , \2205_B[12] , \2210 );
mand \add_15_12/U$16 ( \2397 , \2204_A[12] , \2210 );
mor \add_15_12/U$15 ( \2398 , \2395 , \2396 , \2397 );
mxor \add_15_12/U$13 ( \2399 , \2394 , \2398 );
mbuf \add_15_12/SUM[13] ( \2400_SUM[13] , \2399 );
mand \U$1/U$189 ( \2401 , \2400_SUM[13] , \863 );
mbuf \add_14_12/A[13] ( \2402_A[13] , \a[13] );
mbuf \add_14_12/B[13] ( \2403_B[13] , \c[13] );
mxor \add_14_12/U$14 ( \2404 , \2402_A[13] , \2403_B[13] );
mand \add_14_12/U$18 ( \2405 , \2214_A[12] , \2215_B[12] );
mand \add_14_12/U$17 ( \2406 , \2215_B[12] , \2220 );
mand \add_14_12/U$16 ( \2407 , \2214_A[12] , \2220 );
mor \add_14_12/U$15 ( \2408 , \2405 , \2406 , \2407 );
mxor \add_14_12/U$13 ( \2409 , \2404 , \2408 );
mbuf \add_14_12/SUM[13] ( \2410_SUM[13] , \2409 );
mand \U$1/U$188 ( \2411 , \2410_SUM[13] , \861 );
mand \U$1/U$187 ( \2412 , \d[13] , \859 );
mand \U$1/U$186 ( \2413 , \c[13] , \857 );
mand \U$1/U$185 ( \2414 , \b[13] , \855 );
mand \U$1/U$184 ( \2415 , \a[13] , \853 );
mor \U$1/U$183 ( \2416 , \2229 , \2231 , \2233 , \2235 , \2237 , \2314 , \2391 , \2401 , \2411 , \2412 , \2413 , \2414 , \2415 );
m_DC \n22[14]_g1 ( \2417 , 1'b0 , \876 );
mor \U$5/U$15 ( \2418 , \a[14] , \d[14] );
mand \U$1/U$209 ( \2419 , \2418 , \875 );
mand \U$4/U$15 ( \2420 , \b[14] , \c[14] );
mand \U$1/U$208 ( \2421 , \2420 , \873 );
mor \U$3/U$15 ( \2422 , \a[14] , \b[14] );
mand \U$1/U$207 ( \2423 , \2422 , \871 );
mxor \U$2/U$15 ( \2424 , \c[14] , \d[14] );
mand \U$1/U$206 ( \2425 , \2424 , \869 );
mbuf \mul_17_13/A[14] ( \2426_A[14] , \b[14] );
mand \mul_17_13/U$1394 ( \2427 , \2426_A[14] , \887_B[0] );
mand \mul_17_13/U$1379 ( \2428 , \2238_A[13] , \922_B[1] );
mxor \mul_17_13/U$1314 ( \2429 , \2427 , \2428 );
mand \mul_17_13/U$1318 ( \2430 , \2239 , \2240 );
mand \mul_17_13/U$1317 ( \2431 , \2241 , \2244 );
mor \mul_17_13/U$1315 ( \2432 , \2430 , \2431 );
mxor \mul_17_13/U$1311 ( \2433 , \2429 , \2432 );
mand \mul_17_13/U$1290 ( \2434 , \2062_A[12] , \968_B[2] );
mxor \mul_17_13/U$1229 ( \2435 , \2433 , \2434 );
mand \mul_17_13/U$1233 ( \2436 , \2245 , \2246 );
mand \mul_17_13/U$1232 ( \2437 , \2247 , \2250 );
mor \mul_17_13/U$1230 ( \2438 , \2436 , \2437 );
mxor \mul_17_13/U$1226 ( \2439 , \2435 , \2438 );
mand \mul_17_13/U$1198 ( \2440 , \1898_A[11] , \1030_B[3] );
mxor \mul_17_13/U$1141 ( \2441 , \2439 , \2440 );
mand \mul_17_13/U$1145 ( \2442 , \2251 , \2252 );
mand \mul_17_13/U$1144 ( \2443 , \2253 , \2256 );
mor \mul_17_13/U$1142 ( \2444 , \2442 , \2443 );
mxor \mul_17_13/U$1138 ( \2445 , \2441 , \2444 );
mand \mul_17_13/U$1106 ( \2446 , \1746_A[10] , \1104_B[4] );
mxor \mul_17_13/U$1053 ( \2447 , \2445 , \2446 );
mand \mul_17_13/U$1057 ( \2448 , \2257 , \2258 );
mand \mul_17_13/U$1056 ( \2449 , \2259 , \2262 );
mor \mul_17_13/U$1054 ( \2450 , \2448 , \2449 );
mxor \mul_17_13/U$1050 ( \2451 , \2447 , \2450 );
mand \mul_17_13/U$1014 ( \2452 , \1606_A[9] , \1190_B[5] );
mxor \mul_17_13/U$965 ( \2453 , \2451 , \2452 );
mand \mul_17_13/U$969 ( \2454 , \2263 , \2264 );
mand \mul_17_13/U$968 ( \2455 , \2265 , \2268 );
mor \mul_17_13/U$966 ( \2456 , \2454 , \2455 );
mxor \mul_17_13/U$962 ( \2457 , \2453 , \2456 );
mand \mul_17_13/U$922 ( \2458 , \1478_A[8] , \1288_B[6] );
mxor \mul_17_13/U$877 ( \2459 , \2457 , \2458 );
mand \mul_17_13/U$881 ( \2460 , \2269 , \2270 );
mand \mul_17_13/U$880 ( \2461 , \2271 , \2274 );
mor \mul_17_13/U$878 ( \2462 , \2460 , \2461 );
mxor \mul_17_13/U$874 ( \2463 , \2459 , \2462 );
mand \mul_17_13/U$830 ( \2464 , \1362_A[7] , \1398_B[7] );
mxor \mul_17_13/U$789 ( \2465 , \2463 , \2464 );
mand \mul_17_13/U$793 ( \2466 , \2275 , \2276 );
mand \mul_17_13/U$792 ( \2467 , \2277 , \2280 );
mor \mul_17_13/U$790 ( \2468 , \2466 , \2467 );
mxor \mul_17_13/U$786 ( \2469 , \2465 , \2468 );
mand \mul_17_13/U$738 ( \2470 , \1258_A[6] , \1520_B[8] );
mxor \mul_17_13/U$701 ( \2471 , \2469 , \2470 );
mand \mul_17_13/U$705 ( \2472 , \2281 , \2282 );
mand \mul_17_13/U$704 ( \2473 , \2283 , \2286 );
mor \mul_17_13/U$702 ( \2474 , \2472 , \2473 );
mxor \mul_17_13/U$698 ( \2475 , \2471 , \2474 );
mand \mul_17_13/U$646 ( \2476 , \1166_A[5] , \1654_B[9] );
mxor \mul_17_13/U$613 ( \2477 , \2475 , \2476 );
mand \mul_17_13/U$617 ( \2478 , \2287 , \2288 );
mand \mul_17_13/U$616 ( \2479 , \2289 , \2292 );
mor \mul_17_13/U$614 ( \2480 , \2478 , \2479 );
mxor \mul_17_13/U$610 ( \2481 , \2477 , \2480 );
mand \mul_17_13/U$554 ( \2482 , \1086_A[4] , \1800_B[10] );
mxor \mul_17_13/U$525 ( \2483 , \2481 , \2482 );
mand \mul_17_13/U$529 ( \2484 , \2293 , \2294 );
mand \mul_17_13/U$528 ( \2485 , \2295 , \2298 );
mor \mul_17_13/U$526 ( \2486 , \2484 , \2485 );
mxor \mul_17_13/U$522 ( \2487 , \2483 , \2486 );
mand \mul_17_13/U$462 ( \2488 , \1018_A[3] , \1958_B[11] );
mxor \mul_17_13/U$437 ( \2489 , \2487 , \2488 );
mand \mul_17_13/U$441 ( \2490 , \2299 , \2300 );
mand \mul_17_13/U$440 ( \2491 , \2301 , \2304 );
mor \mul_17_13/U$438 ( \2492 , \2490 , \2491 );
mxor \mul_17_13/U$434 ( \2493 , \2489 , \2492 );
mand \mul_17_13/U$370 ( \2494 , \962_A[2] , \2128_B[12] );
mxor \mul_17_13/U$349 ( \2495 , \2493 , \2494 );
mand \mul_17_13/U$353 ( \2496 , \2305 , \2306 );
mand \mul_17_13/U$352 ( \2497 , \2307 , \2308 );
mor \mul_17_13/U$350 ( \2498 , \2496 , \2497 );
mxor \mul_17_13/U$346 ( \2499 , \2495 , \2498 );
mand \mul_17_13/U$278 ( \2500 , \920_A[1] , \2310_B[13] );
mxor \mul_17_13/U$261 ( \2501 , \2499 , \2500 );
mand \mul_17_13/U$262 ( \2502 , \2309 , \2311 );
mxor \mul_17_13/U$258 ( \2503 , \2501 , \2502 );
mbuf \mul_17_13/B[14] ( \2504_B[14] , \c[14] );
mand \mul_17_13/U$186 ( \2505 , \886_A[0] , \2504_B[14] );
mxor \mul_17_13/U$170 ( \2506 , \2503 , \2505 );
mbuf \mul_17_13/Z[14] ( \2507_Z[14] , \2506 );
mand \U$1/U$205 ( \2508 , \2507_Z[14] , \867 );
mbuf \mul_16_12/A[14] ( \2509_A[14] , \a[14] );
mand \mul_16_12/U$1394 ( \2510 , \2509_A[14] , \892_B[0] );
mand \mul_16_12/U$1379 ( \2511 , \2315_A[13] , \929_B[1] );
mxor \mul_16_12/U$1314 ( \2512 , \2510 , \2511 );
mand \mul_16_12/U$1318 ( \2513 , \2316 , \2317 );
mand \mul_16_12/U$1317 ( \2514 , \2318 , \2321 );
mor \mul_16_12/U$1315 ( \2515 , \2513 , \2514 );
mxor \mul_16_12/U$1311 ( \2516 , \2512 , \2515 );
mand \mul_16_12/U$1290 ( \2517 , \2133_A[12] , \979_B[2] );
mxor \mul_16_12/U$1229 ( \2518 , \2516 , \2517 );
mand \mul_16_12/U$1233 ( \2519 , \2322 , \2323 );
mand \mul_16_12/U$1232 ( \2520 , \2324 , \2327 );
mor \mul_16_12/U$1230 ( \2521 , \2519 , \2520 );
mxor \mul_16_12/U$1226 ( \2522 , \2518 , \2521 );
mand \mul_16_12/U$1198 ( \2523 , \1963_A[11] , \1047_B[3] );
mxor \mul_16_12/U$1141 ( \2524 , \2522 , \2523 );
mand \mul_16_12/U$1145 ( \2525 , \2328 , \2329 );
mand \mul_16_12/U$1144 ( \2526 , \2330 , \2333 );
mor \mul_16_12/U$1142 ( \2527 , \2525 , \2526 );
mxor \mul_16_12/U$1138 ( \2528 , \2524 , \2527 );
mand \mul_16_12/U$1106 ( \2529 , \1805_A[10] , \1127_B[4] );
mxor \mul_16_12/U$1053 ( \2530 , \2528 , \2529 );
mand \mul_16_12/U$1057 ( \2531 , \2334 , \2335 );
mand \mul_16_12/U$1056 ( \2532 , \2336 , \2339 );
mor \mul_16_12/U$1054 ( \2533 , \2531 , \2532 );
mxor \mul_16_12/U$1050 ( \2534 , \2530 , \2533 );
mand \mul_16_12/U$1014 ( \2535 , \1659_A[9] , \1219_B[5] );
mxor \mul_16_12/U$965 ( \2536 , \2534 , \2535 );
mand \mul_16_12/U$969 ( \2537 , \2340 , \2341 );
mand \mul_16_12/U$968 ( \2538 , \2342 , \2345 );
mor \mul_16_12/U$966 ( \2539 , \2537 , \2538 );
mxor \mul_16_12/U$962 ( \2540 , \2536 , \2539 );
mand \mul_16_12/U$922 ( \2541 , \1525_A[8] , \1323_B[6] );
mxor \mul_16_12/U$877 ( \2542 , \2540 , \2541 );
mand \mul_16_12/U$881 ( \2543 , \2346 , \2347 );
mand \mul_16_12/U$880 ( \2544 , \2348 , \2351 );
mor \mul_16_12/U$878 ( \2545 , \2543 , \2544 );
mxor \mul_16_12/U$874 ( \2546 , \2542 , \2545 );
mand \mul_16_12/U$830 ( \2547 , \1403_A[7] , \1439_B[7] );
mxor \mul_16_12/U$789 ( \2548 , \2546 , \2547 );
mand \mul_16_12/U$793 ( \2549 , \2352 , \2353 );
mand \mul_16_12/U$792 ( \2550 , \2354 , \2357 );
mor \mul_16_12/U$790 ( \2551 , \2549 , \2550 );
mxor \mul_16_12/U$786 ( \2552 , \2548 , \2551 );
mand \mul_16_12/U$738 ( \2553 , \1293_A[6] , \1567_B[8] );
mxor \mul_16_12/U$701 ( \2554 , \2552 , \2553 );
mand \mul_16_12/U$705 ( \2555 , \2358 , \2359 );
mand \mul_16_12/U$704 ( \2556 , \2360 , \2363 );
mor \mul_16_12/U$702 ( \2557 , \2555 , \2556 );
mxor \mul_16_12/U$698 ( \2558 , \2554 , \2557 );
mand \mul_16_12/U$646 ( \2559 , \1195_A[5] , \1707_B[9] );
mxor \mul_16_12/U$613 ( \2560 , \2558 , \2559 );
mand \mul_16_12/U$617 ( \2561 , \2364 , \2365 );
mand \mul_16_12/U$616 ( \2562 , \2366 , \2369 );
mor \mul_16_12/U$614 ( \2563 , \2561 , \2562 );
mxor \mul_16_12/U$610 ( \2564 , \2560 , \2563 );
mand \mul_16_12/U$554 ( \2565 , \1109_A[4] , \1859_B[10] );
mxor \mul_16_12/U$525 ( \2566 , \2564 , \2565 );
mand \mul_16_12/U$529 ( \2567 , \2370 , \2371 );
mand \mul_16_12/U$528 ( \2568 , \2372 , \2375 );
mor \mul_16_12/U$526 ( \2569 , \2567 , \2568 );
mxor \mul_16_12/U$522 ( \2570 , \2566 , \2569 );
mand \mul_16_12/U$462 ( \2571 , \1035_A[3] , \2023_B[11] );
mxor \mul_16_12/U$437 ( \2572 , \2570 , \2571 );
mand \mul_16_12/U$441 ( \2573 , \2376 , \2377 );
mand \mul_16_12/U$440 ( \2574 , \2378 , \2381 );
mor \mul_16_12/U$438 ( \2575 , \2573 , \2574 );
mxor \mul_16_12/U$434 ( \2576 , \2572 , \2575 );
mand \mul_16_12/U$370 ( \2577 , \973_A[2] , \2199_B[12] );
mxor \mul_16_12/U$349 ( \2578 , \2576 , \2577 );
mand \mul_16_12/U$353 ( \2579 , \2382 , \2383 );
mand \mul_16_12/U$352 ( \2580 , \2384 , \2385 );
mor \mul_16_12/U$350 ( \2581 , \2579 , \2580 );
mxor \mul_16_12/U$346 ( \2582 , \2578 , \2581 );
mand \mul_16_12/U$278 ( \2583 , \927_A[1] , \2387_B[13] );
mxor \mul_16_12/U$261 ( \2584 , \2582 , \2583 );
mand \mul_16_12/U$262 ( \2585 , \2386 , \2388 );
mxor \mul_16_12/U$258 ( \2586 , \2584 , \2585 );
mbuf \mul_16_12/B[14] ( \2587_B[14] , \d[14] );
mand \mul_16_12/U$186 ( \2588 , \891_A[0] , \2587_B[14] );
mxor \mul_16_12/U$170 ( \2589 , \2586 , \2588 );
mbuf \mul_16_12/Z[14] ( \2590_Z[14] , \2589 );
mand \U$1/U$204 ( \2591 , \2590_Z[14] , \865 );
mbuf \add_15_12/A[14] ( \2592_A[14] , \b[14] );
mbuf \add_15_12/B[14] ( \2593_B[14] , \d[14] );
mxor \add_15_12/U$8 ( \2594 , \2592_A[14] , \2593_B[14] );
mand \add_15_12/U$12 ( \2595 , \2392_A[13] , \2393_B[13] );
mand \add_15_12/U$11 ( \2596 , \2393_B[13] , \2398 );
mand \add_15_12/U$10 ( \2597 , \2392_A[13] , \2398 );
mor \add_15_12/U$9 ( \2598 , \2595 , \2596 , \2597 );
mxor \add_15_12/U$7 ( \2599 , \2594 , \2598 );
mbuf \add_15_12/SUM[14] ( \2600_SUM[14] , \2599 );
mand \U$1/U$203 ( \2601 , \2600_SUM[14] , \863 );
mbuf \add_14_12/A[14] ( \2602_A[14] , \a[14] );
mbuf \add_14_12/B[14] ( \2603_B[14] , \c[14] );
mxor \add_14_12/U$8 ( \2604 , \2602_A[14] , \2603_B[14] );
mand \add_14_12/U$12 ( \2605 , \2402_A[13] , \2403_B[13] );
mand \add_14_12/U$11 ( \2606 , \2403_B[13] , \2408 );
mand \add_14_12/U$10 ( \2607 , \2402_A[13] , \2408 );
mor \add_14_12/U$9 ( \2608 , \2605 , \2606 , \2607 );
mxor \add_14_12/U$7 ( \2609 , \2604 , \2608 );
mbuf \add_14_12/SUM[14] ( \2610_SUM[14] , \2609 );
mand \U$1/U$202 ( \2611 , \2610_SUM[14] , \861 );
mand \U$1/U$201 ( \2612 , \d[14] , \859 );
mand \U$1/U$200 ( \2613 , \c[14] , \857 );
mand \U$1/U$199 ( \2614 , \b[14] , \855 );
mand \U$1/U$198 ( \2615 , \a[14] , \853 );
mor \U$1/U$197 ( \2616 , \2417 , \2419 , \2421 , \2423 , \2425 , \2508 , \2591 , \2601 , \2611 , \2612 , \2613 , \2614 , \2615 );
m_DC \n22[15]_g1 ( \2617 , 1'b0 , \876 );
mor \U$5/U$16 ( \2618 , \a[15] , \d[15] );
mand \U$1/U$223 ( \2619 , \2618 , \875 );
mand \U$4/U$16 ( \2620 , \b[15] , \c[15] );
mand \U$1/U$222 ( \2621 , \2620 , \873 );
mor \U$3/U$16 ( \2622 , \a[15] , \b[15] );
mand \U$1/U$221 ( \2623 , \2622 , \871 );
mxor \U$2/U$16 ( \2624 , \c[15] , \d[15] );
mand \U$1/U$220 ( \2625 , \2624 , \869 );
mbuf \mul_17_13/A[15] ( \2626_A[15] , \b[15] );
mand \mul_17_13/U$1393 ( \2627 , \2626_A[15] , \887_B[0] );
mand \mul_17_13/U$1378 ( \2628 , \2426_A[14] , \922_B[1] );
mxor \mul_17_13/U$1309 ( \2629 , \2627 , \2628 );
mand \mul_17_13/U$1313 ( \2630 , \2427 , \2428 );
mand \mul_17_13/U$1312 ( \2631 , \2429 , \2432 );
mor \mul_17_13/U$1310 ( \2632 , \2630 , \2631 );
mxor \mul_17_13/U$1306 ( \2633 , \2629 , \2632 );
mand \mul_17_13/U$1289 ( \2634 , \2238_A[13] , \968_B[2] );
mxor \mul_17_13/U$1224 ( \2635 , \2633 , \2634 );
mand \mul_17_13/U$1228 ( \2636 , \2433 , \2434 );
mand \mul_17_13/U$1227 ( \2637 , \2435 , \2438 );
mor \mul_17_13/U$1225 ( \2638 , \2636 , \2637 );
mxor \mul_17_13/U$1221 ( \2639 , \2635 , \2638 );
mand \mul_17_13/U$1197 ( \2640 , \2062_A[12] , \1030_B[3] );
mxor \mul_17_13/U$1136 ( \2641 , \2639 , \2640 );
mand \mul_17_13/U$1140 ( \2642 , \2439 , \2440 );
mand \mul_17_13/U$1139 ( \2643 , \2441 , \2444 );
mor \mul_17_13/U$1137 ( \2644 , \2642 , \2643 );
mxor \mul_17_13/U$1133 ( \2645 , \2641 , \2644 );
mand \mul_17_13/U$1105 ( \2646 , \1898_A[11] , \1104_B[4] );
mxor \mul_17_13/U$1048 ( \2647 , \2645 , \2646 );
mand \mul_17_13/U$1052 ( \2648 , \2445 , \2446 );
mand \mul_17_13/U$1051 ( \2649 , \2447 , \2450 );
mor \mul_17_13/U$1049 ( \2650 , \2648 , \2649 );
mxor \mul_17_13/U$1045 ( \2651 , \2647 , \2650 );
mand \mul_17_13/U$1013 ( \2652 , \1746_A[10] , \1190_B[5] );
mxor \mul_17_13/U$960 ( \2653 , \2651 , \2652 );
mand \mul_17_13/U$964 ( \2654 , \2451 , \2452 );
mand \mul_17_13/U$963 ( \2655 , \2453 , \2456 );
mor \mul_17_13/U$961 ( \2656 , \2654 , \2655 );
mxor \mul_17_13/U$957 ( \2657 , \2653 , \2656 );
mand \mul_17_13/U$921 ( \2658 , \1606_A[9] , \1288_B[6] );
mxor \mul_17_13/U$872 ( \2659 , \2657 , \2658 );
mand \mul_17_13/U$876 ( \2660 , \2457 , \2458 );
mand \mul_17_13/U$875 ( \2661 , \2459 , \2462 );
mor \mul_17_13/U$873 ( \2662 , \2660 , \2661 );
mxor \mul_17_13/U$869 ( \2663 , \2659 , \2662 );
mand \mul_17_13/U$829 ( \2664 , \1478_A[8] , \1398_B[7] );
mxor \mul_17_13/U$784 ( \2665 , \2663 , \2664 );
mand \mul_17_13/U$788 ( \2666 , \2463 , \2464 );
mand \mul_17_13/U$787 ( \2667 , \2465 , \2468 );
mor \mul_17_13/U$785 ( \2668 , \2666 , \2667 );
mxor \mul_17_13/U$781 ( \2669 , \2665 , \2668 );
mand \mul_17_13/U$737 ( \2670 , \1362_A[7] , \1520_B[8] );
mxor \mul_17_13/U$696 ( \2671 , \2669 , \2670 );
mand \mul_17_13/U$700 ( \2672 , \2469 , \2470 );
mand \mul_17_13/U$699 ( \2673 , \2471 , \2474 );
mor \mul_17_13/U$697 ( \2674 , \2672 , \2673 );
mxor \mul_17_13/U$693 ( \2675 , \2671 , \2674 );
mand \mul_17_13/U$645 ( \2676 , \1258_A[6] , \1654_B[9] );
mxor \mul_17_13/U$608 ( \2677 , \2675 , \2676 );
mand \mul_17_13/U$612 ( \2678 , \2475 , \2476 );
mand \mul_17_13/U$611 ( \2679 , \2477 , \2480 );
mor \mul_17_13/U$609 ( \2680 , \2678 , \2679 );
mxor \mul_17_13/U$605 ( \2681 , \2677 , \2680 );
mand \mul_17_13/U$553 ( \2682 , \1166_A[5] , \1800_B[10] );
mxor \mul_17_13/U$520 ( \2683 , \2681 , \2682 );
mand \mul_17_13/U$524 ( \2684 , \2481 , \2482 );
mand \mul_17_13/U$523 ( \2685 , \2483 , \2486 );
mor \mul_17_13/U$521 ( \2686 , \2684 , \2685 );
mxor \mul_17_13/U$517 ( \2687 , \2683 , \2686 );
mand \mul_17_13/U$461 ( \2688 , \1086_A[4] , \1958_B[11] );
mxor \mul_17_13/U$432 ( \2689 , \2687 , \2688 );
mand \mul_17_13/U$436 ( \2690 , \2487 , \2488 );
mand \mul_17_13/U$435 ( \2691 , \2489 , \2492 );
mor \mul_17_13/U$433 ( \2692 , \2690 , \2691 );
mxor \mul_17_13/U$429 ( \2693 , \2689 , \2692 );
mand \mul_17_13/U$369 ( \2694 , \1018_A[3] , \2128_B[12] );
mxor \mul_17_13/U$344 ( \2695 , \2693 , \2694 );
mand \mul_17_13/U$348 ( \2696 , \2493 , \2494 );
mand \mul_17_13/U$347 ( \2697 , \2495 , \2498 );
mor \mul_17_13/U$345 ( \2698 , \2696 , \2697 );
mxor \mul_17_13/U$341 ( \2699 , \2695 , \2698 );
mand \mul_17_13/U$277 ( \2700 , \962_A[2] , \2310_B[13] );
mxor \mul_17_13/U$256 ( \2701 , \2699 , \2700 );
mand \mul_17_13/U$260 ( \2702 , \2499 , \2500 );
mand \mul_17_13/U$259 ( \2703 , \2501 , \2502 );
mor \mul_17_13/U$257 ( \2704 , \2702 , \2703 );
mxor \mul_17_13/U$253 ( \2705 , \2701 , \2704 );
mand \mul_17_13/U$185 ( \2706 , \920_A[1] , \2504_B[14] );
mxor \mul_17_13/U$168 ( \2707 , \2705 , \2706 );
mand \mul_17_13/U$169 ( \2708 , \2503 , \2505 );
mxor \mul_17_13/U$165 ( \2709 , \2707 , \2708 );
mbuf \mul_17_13/B[15] ( \2710_B[15] , \c[15] );
mand \mul_17_13/U$93 ( \2711 , \886_A[0] , \2710_B[15] );
mxor \mul_17_13/U$77 ( \2712 , \2709 , \2711 );
mbuf \mul_17_13/Z[15] ( \2713_Z[15] , \2712 );
mand \U$1/U$219 ( \2714 , \2713_Z[15] , \867 );
mbuf \mul_16_12/A[15] ( \2715_A[15] , \a[15] );
mand \mul_16_12/U$1393 ( \2716 , \2715_A[15] , \892_B[0] );
mand \mul_16_12/U$1378 ( \2717 , \2509_A[14] , \929_B[1] );
mxor \mul_16_12/U$1309 ( \2718 , \2716 , \2717 );
mand \mul_16_12/U$1313 ( \2719 , \2510 , \2511 );
mand \mul_16_12/U$1312 ( \2720 , \2512 , \2515 );
mor \mul_16_12/U$1310 ( \2721 , \2719 , \2720 );
mxor \mul_16_12/U$1306 ( \2722 , \2718 , \2721 );
mand \mul_16_12/U$1289 ( \2723 , \2315_A[13] , \979_B[2] );
mxor \mul_16_12/U$1224 ( \2724 , \2722 , \2723 );
mand \mul_16_12/U$1228 ( \2725 , \2516 , \2517 );
mand \mul_16_12/U$1227 ( \2726 , \2518 , \2521 );
mor \mul_16_12/U$1225 ( \2727 , \2725 , \2726 );
mxor \mul_16_12/U$1221 ( \2728 , \2724 , \2727 );
mand \mul_16_12/U$1197 ( \2729 , \2133_A[12] , \1047_B[3] );
mxor \mul_16_12/U$1136 ( \2730 , \2728 , \2729 );
mand \mul_16_12/U$1140 ( \2731 , \2522 , \2523 );
mand \mul_16_12/U$1139 ( \2732 , \2524 , \2527 );
mor \mul_16_12/U$1137 ( \2733 , \2731 , \2732 );
mxor \mul_16_12/U$1133 ( \2734 , \2730 , \2733 );
mand \mul_16_12/U$1105 ( \2735 , \1963_A[11] , \1127_B[4] );
mxor \mul_16_12/U$1048 ( \2736 , \2734 , \2735 );
mand \mul_16_12/U$1052 ( \2737 , \2528 , \2529 );
mand \mul_16_12/U$1051 ( \2738 , \2530 , \2533 );
mor \mul_16_12/U$1049 ( \2739 , \2737 , \2738 );
mxor \mul_16_12/U$1045 ( \2740 , \2736 , \2739 );
mand \mul_16_12/U$1013 ( \2741 , \1805_A[10] , \1219_B[5] );
mxor \mul_16_12/U$960 ( \2742 , \2740 , \2741 );
mand \mul_16_12/U$964 ( \2743 , \2534 , \2535 );
mand \mul_16_12/U$963 ( \2744 , \2536 , \2539 );
mor \mul_16_12/U$961 ( \2745 , \2743 , \2744 );
mxor \mul_16_12/U$957 ( \2746 , \2742 , \2745 );
mand \mul_16_12/U$921 ( \2747 , \1659_A[9] , \1323_B[6] );
mxor \mul_16_12/U$872 ( \2748 , \2746 , \2747 );
mand \mul_16_12/U$876 ( \2749 , \2540 , \2541 );
mand \mul_16_12/U$875 ( \2750 , \2542 , \2545 );
mor \mul_16_12/U$873 ( \2751 , \2749 , \2750 );
mxor \mul_16_12/U$869 ( \2752 , \2748 , \2751 );
mand \mul_16_12/U$829 ( \2753 , \1525_A[8] , \1439_B[7] );
mxor \mul_16_12/U$784 ( \2754 , \2752 , \2753 );
mand \mul_16_12/U$788 ( \2755 , \2546 , \2547 );
mand \mul_16_12/U$787 ( \2756 , \2548 , \2551 );
mor \mul_16_12/U$785 ( \2757 , \2755 , \2756 );
mxor \mul_16_12/U$781 ( \2758 , \2754 , \2757 );
mand \mul_16_12/U$737 ( \2759 , \1403_A[7] , \1567_B[8] );
mxor \mul_16_12/U$696 ( \2760 , \2758 , \2759 );
mand \mul_16_12/U$700 ( \2761 , \2552 , \2553 );
mand \mul_16_12/U$699 ( \2762 , \2554 , \2557 );
mor \mul_16_12/U$697 ( \2763 , \2761 , \2762 );
mxor \mul_16_12/U$693 ( \2764 , \2760 , \2763 );
mand \mul_16_12/U$645 ( \2765 , \1293_A[6] , \1707_B[9] );
mxor \mul_16_12/U$608 ( \2766 , \2764 , \2765 );
mand \mul_16_12/U$612 ( \2767 , \2558 , \2559 );
mand \mul_16_12/U$611 ( \2768 , \2560 , \2563 );
mor \mul_16_12/U$609 ( \2769 , \2767 , \2768 );
mxor \mul_16_12/U$605 ( \2770 , \2766 , \2769 );
mand \mul_16_12/U$553 ( \2771 , \1195_A[5] , \1859_B[10] );
mxor \mul_16_12/U$520 ( \2772 , \2770 , \2771 );
mand \mul_16_12/U$524 ( \2773 , \2564 , \2565 );
mand \mul_16_12/U$523 ( \2774 , \2566 , \2569 );
mor \mul_16_12/U$521 ( \2775 , \2773 , \2774 );
mxor \mul_16_12/U$517 ( \2776 , \2772 , \2775 );
mand \mul_16_12/U$461 ( \2777 , \1109_A[4] , \2023_B[11] );
mxor \mul_16_12/U$432 ( \2778 , \2776 , \2777 );
mand \mul_16_12/U$436 ( \2779 , \2570 , \2571 );
mand \mul_16_12/U$435 ( \2780 , \2572 , \2575 );
mor \mul_16_12/U$433 ( \2781 , \2779 , \2780 );
mxor \mul_16_12/U$429 ( \2782 , \2778 , \2781 );
mand \mul_16_12/U$369 ( \2783 , \1035_A[3] , \2199_B[12] );
mxor \mul_16_12/U$344 ( \2784 , \2782 , \2783 );
mand \mul_16_12/U$348 ( \2785 , \2576 , \2577 );
mand \mul_16_12/U$347 ( \2786 , \2578 , \2581 );
mor \mul_16_12/U$345 ( \2787 , \2785 , \2786 );
mxor \mul_16_12/U$341 ( \2788 , \2784 , \2787 );
mand \mul_16_12/U$277 ( \2789 , \973_A[2] , \2387_B[13] );
mxor \mul_16_12/U$256 ( \2790 , \2788 , \2789 );
mand \mul_16_12/U$260 ( \2791 , \2582 , \2583 );
mand \mul_16_12/U$259 ( \2792 , \2584 , \2585 );
mor \mul_16_12/U$257 ( \2793 , \2791 , \2792 );
mxor \mul_16_12/U$253 ( \2794 , \2790 , \2793 );
mand \mul_16_12/U$185 ( \2795 , \927_A[1] , \2587_B[14] );
mxor \mul_16_12/U$168 ( \2796 , \2794 , \2795 );
mand \mul_16_12/U$169 ( \2797 , \2586 , \2588 );
mxor \mul_16_12/U$165 ( \2798 , \2796 , \2797 );
mbuf \mul_16_12/B[15] ( \2799_B[15] , \d[15] );
mand \mul_16_12/U$93 ( \2800 , \891_A[0] , \2799_B[15] );
mxor \mul_16_12/U$77 ( \2801 , \2798 , \2800 );
mbuf \mul_16_12/Z[15] ( \2802_Z[15] , \2801 );
mand \U$1/U$218 ( \2803 , \2802_Z[15] , \865 );
mbuf \add_15_12/A[15] ( \2804_A[15] , \b[15] );
mbuf \add_15_12/B[15] ( \2805_B[15] , \d[15] );
mxor \add_15_12/U$2 ( \2806 , \2804_A[15] , \2805_B[15] );
mand \add_15_12/U$6 ( \2807 , \2592_A[14] , \2593_B[14] );
mand \add_15_12/U$5 ( \2808 , \2593_B[14] , \2598 );
mand \add_15_12/U$4 ( \2809 , \2592_A[14] , \2598 );
mor \add_15_12/U$3 ( \2810 , \2807 , \2808 , \2809 );
mxor \add_15_12/U$1 ( \2811 , \2806 , \2810 );
mbuf \add_15_12/SUM[15] ( \2812_SUM[15] , \2811 );
mand \U$1/U$217 ( \2813 , \2812_SUM[15] , \863 );
mbuf \add_14_12/A[15] ( \2814_A[15] , \a[15] );
mbuf \add_14_12/B[15] ( \2815_B[15] , \c[15] );
mxor \add_14_12/U$2 ( \2816 , \2814_A[15] , \2815_B[15] );
mand \add_14_12/U$6 ( \2817 , \2602_A[14] , \2603_B[14] );
mand \add_14_12/U$5 ( \2818 , \2603_B[14] , \2608 );
mand \add_14_12/U$4 ( \2819 , \2602_A[14] , \2608 );
mor \add_14_12/U$3 ( \2820 , \2817 , \2818 , \2819 );
mxor \add_14_12/U$1 ( \2821 , \2816 , \2820 );
mbuf \add_14_12/SUM[15] ( \2822_SUM[15] , \2821 );
mand \U$1/U$216 ( \2823 , \2822_SUM[15] , \861 );
mand \U$1/U$215 ( \2824 , \d[15] , \859 );
mand \U$1/U$214 ( \2825 , \c[15] , \857 );
mand \U$1/U$213 ( \2826 , \b[15] , \855 );
mand \U$1/U$212 ( \2827 , \a[15] , \853 );
mor \U$1/U$211 ( \2828 , \2617 , \2619 , \2621 , \2623 , \2625 , \2714 , \2803 , \2813 , \2823 , \2824 , \2825 , \2826 , \2827 );
mbuf \add_7_12/A[15] ( \2829_A[15] , \c[15] );
mbuf \add_7_12/B[15] ( \2830_B[15] , \d[15] );
mand \add_7_12/U$4 ( \2831 , \2829_A[15] , \2830_B[15] );
mbuf \add_7_12/A[14] ( \2832_A[14] , \c[14] );
mbuf \add_7_12/B[14] ( \2833_B[14] , \d[14] );
mand \add_7_12/U$10 ( \2834 , \2832_A[14] , \2833_B[14] );
mbuf \add_7_12/A[13] ( \2835_A[13] , \c[13] );
mbuf \add_7_12/B[13] ( \2836_B[13] , \d[13] );
mand \add_7_12/U$16 ( \2837 , \2835_A[13] , \2836_B[13] );
mbuf \add_7_12/A[12] ( \2838_A[12] , \c[12] );
mbuf \add_7_12/B[12] ( \2839_B[12] , \d[12] );
mand \add_7_12/U$22 ( \2840 , \2838_A[12] , \2839_B[12] );
mbuf \add_7_12/A[11] ( \2841_A[11] , \c[11] );
mbuf \add_7_12/B[11] ( \2842_B[11] , \d[11] );
mand \add_7_12/U$28 ( \2843 , \2841_A[11] , \2842_B[11] );
mbuf \add_7_12/A[10] ( \2844_A[10] , \c[10] );
mbuf \add_7_12/B[10] ( \2845_B[10] , \d[10] );
mand \add_7_12/U$34 ( \2846 , \2844_A[10] , \2845_B[10] );
mbuf \add_7_12/A[9] ( \2847_A[9] , \c[9] );
mbuf \add_7_12/B[9] ( \2848_B[9] , \d[9] );
mand \add_7_12/U$40 ( \2849 , \2847_A[9] , \2848_B[9] );
mbuf \add_7_12/A[8] ( \2850_A[8] , \c[8] );
mbuf \add_7_12/B[8] ( \2851_B[8] , \d[8] );
mand \add_7_12/U$46 ( \2852 , \2850_A[8] , \2851_B[8] );
mbuf \add_7_12/A[7] ( \2853_A[7] , \c[7] );
mbuf \add_7_12/B[7] ( \2854_B[7] , \d[7] );
mand \add_7_12/U$52 ( \2855 , \2853_A[7] , \2854_B[7] );
mbuf \add_7_12/A[6] ( \2856_A[6] , \c[6] );
mbuf \add_7_12/B[6] ( \2857_B[6] , \d[6] );
mand \add_7_12/U$58 ( \2858 , \2856_A[6] , \2857_B[6] );
mbuf \add_7_12/A[5] ( \2859_A[5] , \c[5] );
mbuf \add_7_12/B[5] ( \2860_B[5] , \d[5] );
mand \add_7_12/U$64 ( \2861 , \2859_A[5] , \2860_B[5] );
mbuf \add_7_12/A[4] ( \2862_A[4] , \c[4] );
mbuf \add_7_12/B[4] ( \2863_B[4] , \d[4] );
mand \add_7_12/U$70 ( \2864 , \2862_A[4] , \2863_B[4] );
mbuf \add_7_12/A[3] ( \2865_A[3] , \c[3] );
mbuf \add_7_12/B[3] ( \2866_B[3] , \d[3] );
mand \add_7_12/U$76 ( \2867 , \2865_A[3] , \2866_B[3] );
mbuf \add_7_12/A[2] ( \2868_A[2] , \c[2] );
mbuf \add_7_12/B[2] ( \2869_B[2] , \d[2] );
mand \add_7_12/U$82 ( \2870 , \2868_A[2] , \2869_B[2] );
mbuf \add_7_12/A[1] ( \2871_A[1] , \c[1] );
mbuf \add_7_12/B[1] ( \2872_B[1] , \d[1] );
mand \add_7_12/U$88 ( \2873 , \2871_A[1] , \2872_B[1] );
mbuf \add_7_12/A[0] ( \2874_A[0] , \c[0] );
mbuf \add_7_12/B[0] ( \2875_B[0] , \d[0] );
mand \add_7_12/U$91 ( \2876 , \2874_A[0] , \2875_B[0] );
mand \add_7_12/U$87 ( \2877 , \2872_B[1] , \2876 );
mand \add_7_12/U$86 ( \2878 , \2871_A[1] , \2876 );
mor \add_7_12/U$85 ( \2879 , \2873 , \2877 , \2878 );
mand \add_7_12/U$81 ( \2880 , \2869_B[2] , \2879 );
mand \add_7_12/U$80 ( \2881 , \2868_A[2] , \2879 );
mor \add_7_12/U$79 ( \2882 , \2870 , \2880 , \2881 );
mand \add_7_12/U$75 ( \2883 , \2866_B[3] , \2882 );
mand \add_7_12/U$74 ( \2884 , \2865_A[3] , \2882 );
mor \add_7_12/U$73 ( \2885 , \2867 , \2883 , \2884 );
mand \add_7_12/U$69 ( \2886 , \2863_B[4] , \2885 );
mand \add_7_12/U$68 ( \2887 , \2862_A[4] , \2885 );
mor \add_7_12/U$67 ( \2888 , \2864 , \2886 , \2887 );
mand \add_7_12/U$63 ( \2889 , \2860_B[5] , \2888 );
mand \add_7_12/U$62 ( \2890 , \2859_A[5] , \2888 );
mor \add_7_12/U$61 ( \2891 , \2861 , \2889 , \2890 );
mand \add_7_12/U$57 ( \2892 , \2857_B[6] , \2891 );
mand \add_7_12/U$56 ( \2893 , \2856_A[6] , \2891 );
mor \add_7_12/U$55 ( \2894 , \2858 , \2892 , \2893 );
mand \add_7_12/U$51 ( \2895 , \2854_B[7] , \2894 );
mand \add_7_12/U$50 ( \2896 , \2853_A[7] , \2894 );
mor \add_7_12/U$49 ( \2897 , \2855 , \2895 , \2896 );
mand \add_7_12/U$45 ( \2898 , \2851_B[8] , \2897 );
mand \add_7_12/U$44 ( \2899 , \2850_A[8] , \2897 );
mor \add_7_12/U$43 ( \2900 , \2852 , \2898 , \2899 );
mand \add_7_12/U$39 ( \2901 , \2848_B[9] , \2900 );
mand \add_7_12/U$38 ( \2902 , \2847_A[9] , \2900 );
mor \add_7_12/U$37 ( \2903 , \2849 , \2901 , \2902 );
mand \add_7_12/U$33 ( \2904 , \2845_B[10] , \2903 );
mand \add_7_12/U$32 ( \2905 , \2844_A[10] , \2903 );
mor \add_7_12/U$31 ( \2906 , \2846 , \2904 , \2905 );
mand \add_7_12/U$27 ( \2907 , \2842_B[11] , \2906 );
mand \add_7_12/U$26 ( \2908 , \2841_A[11] , \2906 );
mor \add_7_12/U$25 ( \2909 , \2843 , \2907 , \2908 );
mand \add_7_12/U$21 ( \2910 , \2839_B[12] , \2909 );
mand \add_7_12/U$20 ( \2911 , \2838_A[12] , \2909 );
mor \add_7_12/U$19 ( \2912 , \2840 , \2910 , \2911 );
mand \add_7_12/U$15 ( \2913 , \2836_B[13] , \2912 );
mand \add_7_12/U$14 ( \2914 , \2835_A[13] , \2912 );
mor \add_7_12/U$13 ( \2915 , \2837 , \2913 , \2914 );
mand \add_7_12/U$9 ( \2916 , \2833_B[14] , \2915 );
mand \add_7_12/U$8 ( \2917 , \2832_A[14] , \2915 );
mor \add_7_12/U$7 ( \2918 , \2834 , \2916 , \2917 );
mand \add_7_12/U$3 ( \2919 , \2830_B[15] , \2918 );
mand \add_7_12/U$2 ( \2920 , \2829_A[15] , \2918 );
mor \add_7_12/U$1 ( \2921 , \2831 , \2919 , \2920 );
mbuf \add_7_12/SUM[16] ( \2922_SUM[16] , \2921 );
mbuf \mul_7_15/A[16] ( \2923_A[16] , \2922_SUM[16] );
mxor \add_7_12/U$6 ( \2924 , \2829_A[15] , \2830_B[15] );
mxor \add_7_12/U$5 ( \2925 , \2924 , \2918 );
mbuf \add_7_12/SUM[15] ( \2926_SUM[15] , \2925 );
mbuf \mul_7_15/A[15] ( \2927_A[15] , \2926_SUM[15] );
mxor \add_7_12/U$12 ( \2928 , \2832_A[14] , \2833_B[14] );
mxor \add_7_12/U$11 ( \2929 , \2928 , \2915 );
mbuf \add_7_12/SUM[14] ( \2930_SUM[14] , \2929 );
mbuf \mul_7_15/A[14] ( \2931_A[14] , \2930_SUM[14] );
mxor \add_7_12/U$18 ( \2932 , \2835_A[13] , \2836_B[13] );
mxor \add_7_12/U$17 ( \2933 , \2932 , \2912 );
mbuf \add_7_12/SUM[13] ( \2934_SUM[13] , \2933 );
mbuf \mul_7_15/A[13] ( \2935_A[13] , \2934_SUM[13] );
mxor \add_7_12/U$24 ( \2936 , \2838_A[12] , \2839_B[12] );
mxor \add_7_12/U$23 ( \2937 , \2936 , \2909 );
mbuf \add_7_12/SUM[12] ( \2938_SUM[12] , \2937 );
mbuf \mul_7_15/A[12] ( \2939_A[12] , \2938_SUM[12] );
mxor \add_7_12/U$30 ( \2940 , \2841_A[11] , \2842_B[11] );
mxor \add_7_12/U$29 ( \2941 , \2940 , \2906 );
mbuf \add_7_12/SUM[11] ( \2942_SUM[11] , \2941 );
mbuf \mul_7_15/A[11] ( \2943_A[11] , \2942_SUM[11] );
mxor \add_7_12/U$36 ( \2944 , \2844_A[10] , \2845_B[10] );
mxor \add_7_12/U$35 ( \2945 , \2944 , \2903 );
mbuf \add_7_12/SUM[10] ( \2946_SUM[10] , \2945 );
mbuf \mul_7_15/A[10] ( \2947_A[10] , \2946_SUM[10] );
mxor \add_7_12/U$42 ( \2948 , \2847_A[9] , \2848_B[9] );
mxor \add_7_12/U$41 ( \2949 , \2948 , \2900 );
mbuf \add_7_12/SUM[9] ( \2950_SUM[9] , \2949 );
mbuf \mul_7_15/A[9] ( \2951_A[9] , \2950_SUM[9] );
mxor \add_7_12/U$48 ( \2952 , \2850_A[8] , \2851_B[8] );
mxor \add_7_12/U$47 ( \2953 , \2952 , \2897 );
mbuf \add_7_12/SUM[8] ( \2954_SUM[8] , \2953 );
mbuf \mul_7_15/A[8] ( \2955_A[8] , \2954_SUM[8] );
mxor \add_7_12/U$54 ( \2956 , \2853_A[7] , \2854_B[7] );
mxor \add_7_12/U$53 ( \2957 , \2956 , \2894 );
mbuf \add_7_12/SUM[7] ( \2958_SUM[7] , \2957 );
mbuf \mul_7_15/A[7] ( \2959_A[7] , \2958_SUM[7] );
mxor \add_7_12/U$60 ( \2960 , \2856_A[6] , \2857_B[6] );
mxor \add_7_12/U$59 ( \2961 , \2960 , \2891 );
mbuf \add_7_12/SUM[6] ( \2962_SUM[6] , \2961 );
mbuf \mul_7_15/A[6] ( \2963_A[6] , \2962_SUM[6] );
mxor \add_7_12/U$66 ( \2964 , \2859_A[5] , \2860_B[5] );
mxor \add_7_12/U$65 ( \2965 , \2964 , \2888 );
mbuf \add_7_12/SUM[5] ( \2966_SUM[5] , \2965 );
mbuf \mul_7_15/A[5] ( \2967_A[5] , \2966_SUM[5] );
mxor \add_7_12/U$72 ( \2968 , \2862_A[4] , \2863_B[4] );
mxor \add_7_12/U$71 ( \2969 , \2968 , \2885 );
mbuf \add_7_12/SUM[4] ( \2970_SUM[4] , \2969 );
mbuf \mul_7_15/A[4] ( \2971_A[4] , \2970_SUM[4] );
mxor \add_7_12/U$78 ( \2972 , \2865_A[3] , \2866_B[3] );
mxor \add_7_12/U$77 ( \2973 , \2972 , \2882 );
mbuf \add_7_12/SUM[3] ( \2974_SUM[3] , \2973 );
mbuf \mul_7_15/A[3] ( \2975_A[3] , \2974_SUM[3] );
mxor \add_7_12/U$84 ( \2976 , \2868_A[2] , \2869_B[2] );
mxor \add_7_12/U$83 ( \2977 , \2976 , \2879 );
mbuf \add_7_12/SUM[2] ( \2978_SUM[2] , \2977 );
mbuf \mul_7_15/A[2] ( \2979_A[2] , \2978_SUM[2] );
mxor \add_7_12/U$90 ( \2980 , \2871_A[1] , \2872_B[1] );
mxor \add_7_12/U$89 ( \2981 , \2980 , \2876 );
mbuf \add_7_12/SUM[1] ( \2982_SUM[1] , \2981 );
mbuf \mul_7_15/A[1] ( \2983_A[1] , \2982_SUM[1] );
mxor \add_7_12/U$92 ( \2984 , \2874_A[0] , \2875_B[0] );
mbuf \add_7_12/SUM[0] ( \2985_SUM[0] , \2984 );
mbuf \mul_7_15/A[0] ( \2986_A[0] , \2985_SUM[0] );
mbuf \mul_7_15/B[15] ( \2987_B[15] , \2828 );
mbuf \mul_7_15/B[14] ( \2988_B[14] , \2616 );
mbuf \mul_7_15/B[13] ( \2989_B[13] , \2416 );
mbuf \mul_7_15/B[12] ( \2990_B[12] , \2228 );
mbuf \mul_7_15/B[11] ( \2991_B[11] , \2052 );
mbuf \mul_7_15/B[10] ( \2992_B[10] , \1888 );
mbuf \mul_7_15/B[9] ( \2993_B[9] , \1736 );
mbuf \mul_7_15/B[8] ( \2994_B[8] , \1596 );
mbuf \mul_7_15/B[7] ( \2995_B[7] , \1468 );
mbuf \mul_7_15/B[6] ( \2996_B[6] , \1352 );
mbuf \mul_7_15/B[5] ( \2997_B[5] , \1248 );
mbuf \mul_7_15/B[4] ( \2998_B[4] , \1156 );
mbuf \mul_7_15/B[3] ( \2999_B[3] , \1076 );
mbuf \mul_7_15/B[2] ( \3000_B[2] , \1008 );
mbuf \mul_7_15/B[1] ( \3001_B[1] , \952 );
mbuf \mul_7_15/B[0] ( \3002_B[0] , \910 );
mand \mul_7_15/U$1466 ( \3003 , \2923_A[16] , \3001_B[1] );
mand \mul_7_15/U$1483 ( \3004 , \2923_A[16] , \3002_B[0] );
mand \mul_7_15/U$1467 ( \3005 , \2927_A[15] , \3001_B[1] );
mand \mul_7_15/U$1392 ( \3006 , \3004 , \3005 );
mxor \mul_7_15/U$1393 ( \3007 , \3004 , \3005 );
mand \mul_7_15/U$1484 ( \3008 , \2927_A[15] , \3002_B[0] );
mand \mul_7_15/U$1468 ( \3009 , \2931_A[14] , \3001_B[1] );
mand \mul_7_15/U$1397 ( \3010 , \3008 , \3009 );
mxor \mul_7_15/U$1398 ( \3011 , \3008 , \3009 );
mand \mul_7_15/U$1485 ( \3012 , \2931_A[14] , \3002_B[0] );
mand \mul_7_15/U$1469 ( \3013 , \2935_A[13] , \3001_B[1] );
mand \mul_7_15/U$1402 ( \3014 , \3012 , \3013 );
mxor \mul_7_15/U$1403 ( \3015 , \3012 , \3013 );
mand \mul_7_15/U$1486 ( \3016 , \2935_A[13] , \3002_B[0] );
mand \mul_7_15/U$1470 ( \3017 , \2939_A[12] , \3001_B[1] );
mand \mul_7_15/U$1407 ( \3018 , \3016 , \3017 );
mxor \mul_7_15/U$1408 ( \3019 , \3016 , \3017 );
mand \mul_7_15/U$1487 ( \3020 , \2939_A[12] , \3002_B[0] );
mand \mul_7_15/U$1471 ( \3021 , \2943_A[11] , \3001_B[1] );
mand \mul_7_15/U$1412 ( \3022 , \3020 , \3021 );
mxor \mul_7_15/U$1413 ( \3023 , \3020 , \3021 );
mand \mul_7_15/U$1488 ( \3024 , \2943_A[11] , \3002_B[0] );
mand \mul_7_15/U$1472 ( \3025 , \2947_A[10] , \3001_B[1] );
mand \mul_7_15/U$1417 ( \3026 , \3024 , \3025 );
mxor \mul_7_15/U$1418 ( \3027 , \3024 , \3025 );
mand \mul_7_15/U$1489 ( \3028 , \2947_A[10] , \3002_B[0] );
mand \mul_7_15/U$1473 ( \3029 , \2951_A[9] , \3001_B[1] );
mand \mul_7_15/U$1422 ( \3030 , \3028 , \3029 );
mxor \mul_7_15/U$1423 ( \3031 , \3028 , \3029 );
mand \mul_7_15/U$1490 ( \3032 , \2951_A[9] , \3002_B[0] );
mand \mul_7_15/U$1474 ( \3033 , \2955_A[8] , \3001_B[1] );
mand \mul_7_15/U$1427 ( \3034 , \3032 , \3033 );
mxor \mul_7_15/U$1428 ( \3035 , \3032 , \3033 );
mand \mul_7_15/U$1491 ( \3036 , \2955_A[8] , \3002_B[0] );
mand \mul_7_15/U$1475 ( \3037 , \2959_A[7] , \3001_B[1] );
mand \mul_7_15/U$1432 ( \3038 , \3036 , \3037 );
mxor \mul_7_15/U$1433 ( \3039 , \3036 , \3037 );
mand \mul_7_15/U$1492 ( \3040 , \2959_A[7] , \3002_B[0] );
mand \mul_7_15/U$1476 ( \3041 , \2963_A[6] , \3001_B[1] );
mand \mul_7_15/U$1437 ( \3042 , \3040 , \3041 );
mxor \mul_7_15/U$1438 ( \3043 , \3040 , \3041 );
mand \mul_7_15/U$1493 ( \3044 , \2963_A[6] , \3002_B[0] );
mand \mul_7_15/U$1477 ( \3045 , \2967_A[5] , \3001_B[1] );
mand \mul_7_15/U$1442 ( \3046 , \3044 , \3045 );
mxor \mul_7_15/U$1443 ( \3047 , \3044 , \3045 );
mand \mul_7_15/U$1494 ( \3048 , \2967_A[5] , \3002_B[0] );
mand \mul_7_15/U$1478 ( \3049 , \2971_A[4] , \3001_B[1] );
mand \mul_7_15/U$1447 ( \3050 , \3048 , \3049 );
mxor \mul_7_15/U$1448 ( \3051 , \3048 , \3049 );
mand \mul_7_15/U$1495 ( \3052 , \2971_A[4] , \3002_B[0] );
mand \mul_7_15/U$1479 ( \3053 , \2975_A[3] , \3001_B[1] );
mand \mul_7_15/U$1452 ( \3054 , \3052 , \3053 );
mxor \mul_7_15/U$1453 ( \3055 , \3052 , \3053 );
mand \mul_7_15/U$1496 ( \3056 , \2975_A[3] , \3002_B[0] );
mand \mul_7_15/U$1480 ( \3057 , \2979_A[2] , \3001_B[1] );
mand \mul_7_15/U$1457 ( \3058 , \3056 , \3057 );
mxor \mul_7_15/U$1458 ( \3059 , \3056 , \3057 );
mand \mul_7_15/U$1497 ( \3060 , \2979_A[2] , \3002_B[0] );
mand \mul_7_15/U$1481 ( \3061 , \2983_A[1] , \3001_B[1] );
mand \mul_7_15/U$1462 ( \3062 , \3060 , \3061 );
mxor \mul_7_15/U$1463 ( \3063 , \3060 , \3061 );
mand \mul_7_15/U$1498 ( \3064 , \2983_A[1] , \3002_B[0] );
mand \mul_7_15/U$1482 ( \3065 , \2986_A[0] , \3001_B[1] );
mand \mul_7_15/U$1464 ( \3066 , \3064 , \3065 );
mand \mul_7_15/U$1461 ( \3067 , \3063 , \3066 );
mor \mul_7_15/U$1459 ( \3068 , \3062 , \3067 );
mand \mul_7_15/U$1456 ( \3069 , \3059 , \3068 );
mor \mul_7_15/U$1454 ( \3070 , \3058 , \3069 );
mand \mul_7_15/U$1451 ( \3071 , \3055 , \3070 );
mor \mul_7_15/U$1449 ( \3072 , \3054 , \3071 );
mand \mul_7_15/U$1446 ( \3073 , \3051 , \3072 );
mor \mul_7_15/U$1444 ( \3074 , \3050 , \3073 );
mand \mul_7_15/U$1441 ( \3075 , \3047 , \3074 );
mor \mul_7_15/U$1439 ( \3076 , \3046 , \3075 );
mand \mul_7_15/U$1436 ( \3077 , \3043 , \3076 );
mor \mul_7_15/U$1434 ( \3078 , \3042 , \3077 );
mand \mul_7_15/U$1431 ( \3079 , \3039 , \3078 );
mor \mul_7_15/U$1429 ( \3080 , \3038 , \3079 );
mand \mul_7_15/U$1426 ( \3081 , \3035 , \3080 );
mor \mul_7_15/U$1424 ( \3082 , \3034 , \3081 );
mand \mul_7_15/U$1421 ( \3083 , \3031 , \3082 );
mor \mul_7_15/U$1419 ( \3084 , \3030 , \3083 );
mand \mul_7_15/U$1416 ( \3085 , \3027 , \3084 );
mor \mul_7_15/U$1414 ( \3086 , \3026 , \3085 );
mand \mul_7_15/U$1411 ( \3087 , \3023 , \3086 );
mor \mul_7_15/U$1409 ( \3088 , \3022 , \3087 );
mand \mul_7_15/U$1406 ( \3089 , \3019 , \3088 );
mor \mul_7_15/U$1404 ( \3090 , \3018 , \3089 );
mand \mul_7_15/U$1401 ( \3091 , \3015 , \3090 );
mor \mul_7_15/U$1399 ( \3092 , \3014 , \3091 );
mand \mul_7_15/U$1396 ( \3093 , \3011 , \3092 );
mor \mul_7_15/U$1394 ( \3094 , \3010 , \3093 );
mand \mul_7_15/U$1391 ( \3095 , \3007 , \3094 );
mor \mul_7_15/U$1389 ( \3096 , \3006 , \3095 );
mand \mul_7_15/U$1388 ( \3097 , \3003 , \3096 );
mand \mul_7_15/U$1370 ( \3098 , \2923_A[16] , \3000_B[2] );
mand \mul_7_15/U$1291 ( \3099 , \3097 , \3098 );
mxor \mul_7_15/U$1292 ( \3100 , \3097 , \3098 );
mxor \mul_7_15/U$1387 ( \3101 , \3003 , \3096 );
mand \mul_7_15/U$1371 ( \3102 , \2927_A[15] , \3000_B[2] );
mand \mul_7_15/U$1296 ( \3103 , \3101 , \3102 );
mxor \mul_7_15/U$1297 ( \3104 , \3101 , \3102 );
mxor \mul_7_15/U$1390 ( \3105 , \3007 , \3094 );
mand \mul_7_15/U$1372 ( \3106 , \2931_A[14] , \3000_B[2] );
mand \mul_7_15/U$1301 ( \3107 , \3105 , \3106 );
mxor \mul_7_15/U$1302 ( \3108 , \3105 , \3106 );
mxor \mul_7_15/U$1395 ( \3109 , \3011 , \3092 );
mand \mul_7_15/U$1373 ( \3110 , \2935_A[13] , \3000_B[2] );
mand \mul_7_15/U$1306 ( \3111 , \3109 , \3110 );
mxor \mul_7_15/U$1307 ( \3112 , \3109 , \3110 );
mxor \mul_7_15/U$1400 ( \3113 , \3015 , \3090 );
mand \mul_7_15/U$1374 ( \3114 , \2939_A[12] , \3000_B[2] );
mand \mul_7_15/U$1311 ( \3115 , \3113 , \3114 );
mxor \mul_7_15/U$1312 ( \3116 , \3113 , \3114 );
mxor \mul_7_15/U$1405 ( \3117 , \3019 , \3088 );
mand \mul_7_15/U$1375 ( \3118 , \2943_A[11] , \3000_B[2] );
mand \mul_7_15/U$1316 ( \3119 , \3117 , \3118 );
mxor \mul_7_15/U$1317 ( \3120 , \3117 , \3118 );
mxor \mul_7_15/U$1410 ( \3121 , \3023 , \3086 );
mand \mul_7_15/U$1376 ( \3122 , \2947_A[10] , \3000_B[2] );
mand \mul_7_15/U$1321 ( \3123 , \3121 , \3122 );
mxor \mul_7_15/U$1322 ( \3124 , \3121 , \3122 );
mxor \mul_7_15/U$1415 ( \3125 , \3027 , \3084 );
mand \mul_7_15/U$1377 ( \3126 , \2951_A[9] , \3000_B[2] );
mand \mul_7_15/U$1326 ( \3127 , \3125 , \3126 );
mxor \mul_7_15/U$1327 ( \3128 , \3125 , \3126 );
mxor \mul_7_15/U$1420 ( \3129 , \3031 , \3082 );
mand \mul_7_15/U$1378 ( \3130 , \2955_A[8] , \3000_B[2] );
mand \mul_7_15/U$1331 ( \3131 , \3129 , \3130 );
mxor \mul_7_15/U$1332 ( \3132 , \3129 , \3130 );
mxor \mul_7_15/U$1425 ( \3133 , \3035 , \3080 );
mand \mul_7_15/U$1379 ( \3134 , \2959_A[7] , \3000_B[2] );
mand \mul_7_15/U$1336 ( \3135 , \3133 , \3134 );
mxor \mul_7_15/U$1337 ( \3136 , \3133 , \3134 );
mxor \mul_7_15/U$1430 ( \3137 , \3039 , \3078 );
mand \mul_7_15/U$1380 ( \3138 , \2963_A[6] , \3000_B[2] );
mand \mul_7_15/U$1341 ( \3139 , \3137 , \3138 );
mxor \mul_7_15/U$1342 ( \3140 , \3137 , \3138 );
mxor \mul_7_15/U$1435 ( \3141 , \3043 , \3076 );
mand \mul_7_15/U$1381 ( \3142 , \2967_A[5] , \3000_B[2] );
mand \mul_7_15/U$1346 ( \3143 , \3141 , \3142 );
mxor \mul_7_15/U$1347 ( \3144 , \3141 , \3142 );
mxor \mul_7_15/U$1440 ( \3145 , \3047 , \3074 );
mand \mul_7_15/U$1382 ( \3146 , \2971_A[4] , \3000_B[2] );
mand \mul_7_15/U$1351 ( \3147 , \3145 , \3146 );
mxor \mul_7_15/U$1352 ( \3148 , \3145 , \3146 );
mxor \mul_7_15/U$1445 ( \3149 , \3051 , \3072 );
mand \mul_7_15/U$1383 ( \3150 , \2975_A[3] , \3000_B[2] );
mand \mul_7_15/U$1356 ( \3151 , \3149 , \3150 );
mxor \mul_7_15/U$1357 ( \3152 , \3149 , \3150 );
mxor \mul_7_15/U$1450 ( \3153 , \3055 , \3070 );
mand \mul_7_15/U$1384 ( \3154 , \2979_A[2] , \3000_B[2] );
mand \mul_7_15/U$1361 ( \3155 , \3153 , \3154 );
mxor \mul_7_15/U$1362 ( \3156 , \3153 , \3154 );
mxor \mul_7_15/U$1455 ( \3157 , \3059 , \3068 );
mand \mul_7_15/U$1385 ( \3158 , \2983_A[1] , \3000_B[2] );
mand \mul_7_15/U$1366 ( \3159 , \3157 , \3158 );
mxor \mul_7_15/U$1367 ( \3160 , \3157 , \3158 );
mxor \mul_7_15/U$1460 ( \3161 , \3063 , \3066 );
mand \mul_7_15/U$1386 ( \3162 , \2986_A[0] , \3000_B[2] );
mand \mul_7_15/U$1368 ( \3163 , \3161 , \3162 );
mand \mul_7_15/U$1365 ( \3164 , \3160 , \3163 );
mor \mul_7_15/U$1363 ( \3165 , \3159 , \3164 );
mand \mul_7_15/U$1360 ( \3166 , \3156 , \3165 );
mor \mul_7_15/U$1358 ( \3167 , \3155 , \3166 );
mand \mul_7_15/U$1355 ( \3168 , \3152 , \3167 );
mor \mul_7_15/U$1353 ( \3169 , \3151 , \3168 );
mand \mul_7_15/U$1350 ( \3170 , \3148 , \3169 );
mor \mul_7_15/U$1348 ( \3171 , \3147 , \3170 );
mand \mul_7_15/U$1345 ( \3172 , \3144 , \3171 );
mor \mul_7_15/U$1343 ( \3173 , \3143 , \3172 );
mand \mul_7_15/U$1340 ( \3174 , \3140 , \3173 );
mor \mul_7_15/U$1338 ( \3175 , \3139 , \3174 );
mand \mul_7_15/U$1335 ( \3176 , \3136 , \3175 );
mor \mul_7_15/U$1333 ( \3177 , \3135 , \3176 );
mand \mul_7_15/U$1330 ( \3178 , \3132 , \3177 );
mor \mul_7_15/U$1328 ( \3179 , \3131 , \3178 );
mand \mul_7_15/U$1325 ( \3180 , \3128 , \3179 );
mor \mul_7_15/U$1323 ( \3181 , \3127 , \3180 );
mand \mul_7_15/U$1320 ( \3182 , \3124 , \3181 );
mor \mul_7_15/U$1318 ( \3183 , \3123 , \3182 );
mand \mul_7_15/U$1315 ( \3184 , \3120 , \3183 );
mor \mul_7_15/U$1313 ( \3185 , \3119 , \3184 );
mand \mul_7_15/U$1310 ( \3186 , \3116 , \3185 );
mor \mul_7_15/U$1308 ( \3187 , \3115 , \3186 );
mand \mul_7_15/U$1305 ( \3188 , \3112 , \3187 );
mor \mul_7_15/U$1303 ( \3189 , \3111 , \3188 );
mand \mul_7_15/U$1300 ( \3190 , \3108 , \3189 );
mor \mul_7_15/U$1298 ( \3191 , \3107 , \3190 );
mand \mul_7_15/U$1295 ( \3192 , \3104 , \3191 );
mor \mul_7_15/U$1293 ( \3193 , \3103 , \3192 );
mand \mul_7_15/U$1290 ( \3194 , \3100 , \3193 );
mor \mul_7_15/U$1288 ( \3195 , \3099 , \3194 );
mand \mul_7_15/U$1271 ( \3196 , \2923_A[16] , \2999_B[3] );
mand \mul_7_15/U$1192 ( \3197 , \3195 , \3196 );
mxor \mul_7_15/U$1193 ( \3198 , \3195 , \3196 );
mxor \mul_7_15/U$1289 ( \3199 , \3100 , \3193 );
mand \mul_7_15/U$1272 ( \3200 , \2927_A[15] , \2999_B[3] );
mand \mul_7_15/U$1197 ( \3201 , \3199 , \3200 );
mxor \mul_7_15/U$1198 ( \3202 , \3199 , \3200 );
mxor \mul_7_15/U$1294 ( \3203 , \3104 , \3191 );
mand \mul_7_15/U$1273 ( \3204 , \2931_A[14] , \2999_B[3] );
mand \mul_7_15/U$1202 ( \3205 , \3203 , \3204 );
mxor \mul_7_15/U$1203 ( \3206 , \3203 , \3204 );
mxor \mul_7_15/U$1299 ( \3207 , \3108 , \3189 );
mand \mul_7_15/U$1274 ( \3208 , \2935_A[13] , \2999_B[3] );
mand \mul_7_15/U$1207 ( \3209 , \3207 , \3208 );
mxor \mul_7_15/U$1208 ( \3210 , \3207 , \3208 );
mxor \mul_7_15/U$1304 ( \3211 , \3112 , \3187 );
mand \mul_7_15/U$1275 ( \3212 , \2939_A[12] , \2999_B[3] );
mand \mul_7_15/U$1212 ( \3213 , \3211 , \3212 );
mxor \mul_7_15/U$1213 ( \3214 , \3211 , \3212 );
mxor \mul_7_15/U$1309 ( \3215 , \3116 , \3185 );
mand \mul_7_15/U$1276 ( \3216 , \2943_A[11] , \2999_B[3] );
mand \mul_7_15/U$1217 ( \3217 , \3215 , \3216 );
mxor \mul_7_15/U$1218 ( \3218 , \3215 , \3216 );
mxor \mul_7_15/U$1314 ( \3219 , \3120 , \3183 );
mand \mul_7_15/U$1277 ( \3220 , \2947_A[10] , \2999_B[3] );
mand \mul_7_15/U$1222 ( \3221 , \3219 , \3220 );
mxor \mul_7_15/U$1223 ( \3222 , \3219 , \3220 );
mxor \mul_7_15/U$1319 ( \3223 , \3124 , \3181 );
mand \mul_7_15/U$1278 ( \3224 , \2951_A[9] , \2999_B[3] );
mand \mul_7_15/U$1227 ( \3225 , \3223 , \3224 );
mxor \mul_7_15/U$1228 ( \3226 , \3223 , \3224 );
mxor \mul_7_15/U$1324 ( \3227 , \3128 , \3179 );
mand \mul_7_15/U$1279 ( \3228 , \2955_A[8] , \2999_B[3] );
mand \mul_7_15/U$1232 ( \3229 , \3227 , \3228 );
mxor \mul_7_15/U$1233 ( \3230 , \3227 , \3228 );
mxor \mul_7_15/U$1329 ( \3231 , \3132 , \3177 );
mand \mul_7_15/U$1280 ( \3232 , \2959_A[7] , \2999_B[3] );
mand \mul_7_15/U$1237 ( \3233 , \3231 , \3232 );
mxor \mul_7_15/U$1238 ( \3234 , \3231 , \3232 );
mxor \mul_7_15/U$1334 ( \3235 , \3136 , \3175 );
mand \mul_7_15/U$1281 ( \3236 , \2963_A[6] , \2999_B[3] );
mand \mul_7_15/U$1242 ( \3237 , \3235 , \3236 );
mxor \mul_7_15/U$1243 ( \3238 , \3235 , \3236 );
mxor \mul_7_15/U$1339 ( \3239 , \3140 , \3173 );
mand \mul_7_15/U$1282 ( \3240 , \2967_A[5] , \2999_B[3] );
mand \mul_7_15/U$1247 ( \3241 , \3239 , \3240 );
mxor \mul_7_15/U$1248 ( \3242 , \3239 , \3240 );
mxor \mul_7_15/U$1344 ( \3243 , \3144 , \3171 );
mand \mul_7_15/U$1283 ( \3244 , \2971_A[4] , \2999_B[3] );
mand \mul_7_15/U$1252 ( \3245 , \3243 , \3244 );
mxor \mul_7_15/U$1253 ( \3246 , \3243 , \3244 );
mxor \mul_7_15/U$1349 ( \3247 , \3148 , \3169 );
mand \mul_7_15/U$1284 ( \3248 , \2975_A[3] , \2999_B[3] );
mand \mul_7_15/U$1257 ( \3249 , \3247 , \3248 );
mxor \mul_7_15/U$1258 ( \3250 , \3247 , \3248 );
mxor \mul_7_15/U$1354 ( \3251 , \3152 , \3167 );
mand \mul_7_15/U$1285 ( \3252 , \2979_A[2] , \2999_B[3] );
mand \mul_7_15/U$1262 ( \3253 , \3251 , \3252 );
mxor \mul_7_15/U$1263 ( \3254 , \3251 , \3252 );
mxor \mul_7_15/U$1359 ( \3255 , \3156 , \3165 );
mand \mul_7_15/U$1286 ( \3256 , \2983_A[1] , \2999_B[3] );
mand \mul_7_15/U$1267 ( \3257 , \3255 , \3256 );
mxor \mul_7_15/U$1268 ( \3258 , \3255 , \3256 );
mxor \mul_7_15/U$1364 ( \3259 , \3160 , \3163 );
mand \mul_7_15/U$1287 ( \3260 , \2986_A[0] , \2999_B[3] );
mand \mul_7_15/U$1269 ( \3261 , \3259 , \3260 );
mand \mul_7_15/U$1266 ( \3262 , \3258 , \3261 );
mor \mul_7_15/U$1264 ( \3263 , \3257 , \3262 );
mand \mul_7_15/U$1261 ( \3264 , \3254 , \3263 );
mor \mul_7_15/U$1259 ( \3265 , \3253 , \3264 );
mand \mul_7_15/U$1256 ( \3266 , \3250 , \3265 );
mor \mul_7_15/U$1254 ( \3267 , \3249 , \3266 );
mand \mul_7_15/U$1251 ( \3268 , \3246 , \3267 );
mor \mul_7_15/U$1249 ( \3269 , \3245 , \3268 );
mand \mul_7_15/U$1246 ( \3270 , \3242 , \3269 );
mor \mul_7_15/U$1244 ( \3271 , \3241 , \3270 );
mand \mul_7_15/U$1241 ( \3272 , \3238 , \3271 );
mor \mul_7_15/U$1239 ( \3273 , \3237 , \3272 );
mand \mul_7_15/U$1236 ( \3274 , \3234 , \3273 );
mor \mul_7_15/U$1234 ( \3275 , \3233 , \3274 );
mand \mul_7_15/U$1231 ( \3276 , \3230 , \3275 );
mor \mul_7_15/U$1229 ( \3277 , \3229 , \3276 );
mand \mul_7_15/U$1226 ( \3278 , \3226 , \3277 );
mor \mul_7_15/U$1224 ( \3279 , \3225 , \3278 );
mand \mul_7_15/U$1221 ( \3280 , \3222 , \3279 );
mor \mul_7_15/U$1219 ( \3281 , \3221 , \3280 );
mand \mul_7_15/U$1216 ( \3282 , \3218 , \3281 );
mor \mul_7_15/U$1214 ( \3283 , \3217 , \3282 );
mand \mul_7_15/U$1211 ( \3284 , \3214 , \3283 );
mor \mul_7_15/U$1209 ( \3285 , \3213 , \3284 );
mand \mul_7_15/U$1206 ( \3286 , \3210 , \3285 );
mor \mul_7_15/U$1204 ( \3287 , \3209 , \3286 );
mand \mul_7_15/U$1201 ( \3288 , \3206 , \3287 );
mor \mul_7_15/U$1199 ( \3289 , \3205 , \3288 );
mand \mul_7_15/U$1196 ( \3290 , \3202 , \3289 );
mor \mul_7_15/U$1194 ( \3291 , \3201 , \3290 );
mand \mul_7_15/U$1191 ( \3292 , \3198 , \3291 );
mor \mul_7_15/U$1189 ( \3293 , \3197 , \3292 );
mand \mul_7_15/U$1172 ( \3294 , \2923_A[16] , \2998_B[4] );
mand \mul_7_15/U$1093 ( \3295 , \3293 , \3294 );
mxor \mul_7_15/U$1094 ( \3296 , \3293 , \3294 );
mxor \mul_7_15/U$1190 ( \3297 , \3198 , \3291 );
mand \mul_7_15/U$1173 ( \3298 , \2927_A[15] , \2998_B[4] );
mand \mul_7_15/U$1098 ( \3299 , \3297 , \3298 );
mxor \mul_7_15/U$1099 ( \3300 , \3297 , \3298 );
mxor \mul_7_15/U$1195 ( \3301 , \3202 , \3289 );
mand \mul_7_15/U$1174 ( \3302 , \2931_A[14] , \2998_B[4] );
mand \mul_7_15/U$1103 ( \3303 , \3301 , \3302 );
mxor \mul_7_15/U$1104 ( \3304 , \3301 , \3302 );
mxor \mul_7_15/U$1200 ( \3305 , \3206 , \3287 );
mand \mul_7_15/U$1175 ( \3306 , \2935_A[13] , \2998_B[4] );
mand \mul_7_15/U$1108 ( \3307 , \3305 , \3306 );
mxor \mul_7_15/U$1109 ( \3308 , \3305 , \3306 );
mxor \mul_7_15/U$1205 ( \3309 , \3210 , \3285 );
mand \mul_7_15/U$1176 ( \3310 , \2939_A[12] , \2998_B[4] );
mand \mul_7_15/U$1113 ( \3311 , \3309 , \3310 );
mxor \mul_7_15/U$1114 ( \3312 , \3309 , \3310 );
mxor \mul_7_15/U$1210 ( \3313 , \3214 , \3283 );
mand \mul_7_15/U$1177 ( \3314 , \2943_A[11] , \2998_B[4] );
mand \mul_7_15/U$1118 ( \3315 , \3313 , \3314 );
mxor \mul_7_15/U$1119 ( \3316 , \3313 , \3314 );
mxor \mul_7_15/U$1215 ( \3317 , \3218 , \3281 );
mand \mul_7_15/U$1178 ( \3318 , \2947_A[10] , \2998_B[4] );
mand \mul_7_15/U$1123 ( \3319 , \3317 , \3318 );
mxor \mul_7_15/U$1124 ( \3320 , \3317 , \3318 );
mxor \mul_7_15/U$1220 ( \3321 , \3222 , \3279 );
mand \mul_7_15/U$1179 ( \3322 , \2951_A[9] , \2998_B[4] );
mand \mul_7_15/U$1128 ( \3323 , \3321 , \3322 );
mxor \mul_7_15/U$1129 ( \3324 , \3321 , \3322 );
mxor \mul_7_15/U$1225 ( \3325 , \3226 , \3277 );
mand \mul_7_15/U$1180 ( \3326 , \2955_A[8] , \2998_B[4] );
mand \mul_7_15/U$1133 ( \3327 , \3325 , \3326 );
mxor \mul_7_15/U$1134 ( \3328 , \3325 , \3326 );
mxor \mul_7_15/U$1230 ( \3329 , \3230 , \3275 );
mand \mul_7_15/U$1181 ( \3330 , \2959_A[7] , \2998_B[4] );
mand \mul_7_15/U$1138 ( \3331 , \3329 , \3330 );
mxor \mul_7_15/U$1139 ( \3332 , \3329 , \3330 );
mxor \mul_7_15/U$1235 ( \3333 , \3234 , \3273 );
mand \mul_7_15/U$1182 ( \3334 , \2963_A[6] , \2998_B[4] );
mand \mul_7_15/U$1143 ( \3335 , \3333 , \3334 );
mxor \mul_7_15/U$1144 ( \3336 , \3333 , \3334 );
mxor \mul_7_15/U$1240 ( \3337 , \3238 , \3271 );
mand \mul_7_15/U$1183 ( \3338 , \2967_A[5] , \2998_B[4] );
mand \mul_7_15/U$1148 ( \3339 , \3337 , \3338 );
mxor \mul_7_15/U$1149 ( \3340 , \3337 , \3338 );
mxor \mul_7_15/U$1245 ( \3341 , \3242 , \3269 );
mand \mul_7_15/U$1184 ( \3342 , \2971_A[4] , \2998_B[4] );
mand \mul_7_15/U$1153 ( \3343 , \3341 , \3342 );
mxor \mul_7_15/U$1154 ( \3344 , \3341 , \3342 );
mxor \mul_7_15/U$1250 ( \3345 , \3246 , \3267 );
mand \mul_7_15/U$1185 ( \3346 , \2975_A[3] , \2998_B[4] );
mand \mul_7_15/U$1158 ( \3347 , \3345 , \3346 );
mxor \mul_7_15/U$1159 ( \3348 , \3345 , \3346 );
mxor \mul_7_15/U$1255 ( \3349 , \3250 , \3265 );
mand \mul_7_15/U$1186 ( \3350 , \2979_A[2] , \2998_B[4] );
mand \mul_7_15/U$1163 ( \3351 , \3349 , \3350 );
mxor \mul_7_15/U$1164 ( \3352 , \3349 , \3350 );
mxor \mul_7_15/U$1260 ( \3353 , \3254 , \3263 );
mand \mul_7_15/U$1187 ( \3354 , \2983_A[1] , \2998_B[4] );
mand \mul_7_15/U$1168 ( \3355 , \3353 , \3354 );
mxor \mul_7_15/U$1169 ( \3356 , \3353 , \3354 );
mxor \mul_7_15/U$1265 ( \3357 , \3258 , \3261 );
mand \mul_7_15/U$1188 ( \3358 , \2986_A[0] , \2998_B[4] );
mand \mul_7_15/U$1170 ( \3359 , \3357 , \3358 );
mand \mul_7_15/U$1167 ( \3360 , \3356 , \3359 );
mor \mul_7_15/U$1165 ( \3361 , \3355 , \3360 );
mand \mul_7_15/U$1162 ( \3362 , \3352 , \3361 );
mor \mul_7_15/U$1160 ( \3363 , \3351 , \3362 );
mand \mul_7_15/U$1157 ( \3364 , \3348 , \3363 );
mor \mul_7_15/U$1155 ( \3365 , \3347 , \3364 );
mand \mul_7_15/U$1152 ( \3366 , \3344 , \3365 );
mor \mul_7_15/U$1150 ( \3367 , \3343 , \3366 );
mand \mul_7_15/U$1147 ( \3368 , \3340 , \3367 );
mor \mul_7_15/U$1145 ( \3369 , \3339 , \3368 );
mand \mul_7_15/U$1142 ( \3370 , \3336 , \3369 );
mor \mul_7_15/U$1140 ( \3371 , \3335 , \3370 );
mand \mul_7_15/U$1137 ( \3372 , \3332 , \3371 );
mor \mul_7_15/U$1135 ( \3373 , \3331 , \3372 );
mand \mul_7_15/U$1132 ( \3374 , \3328 , \3373 );
mor \mul_7_15/U$1130 ( \3375 , \3327 , \3374 );
mand \mul_7_15/U$1127 ( \3376 , \3324 , \3375 );
mor \mul_7_15/U$1125 ( \3377 , \3323 , \3376 );
mand \mul_7_15/U$1122 ( \3378 , \3320 , \3377 );
mor \mul_7_15/U$1120 ( \3379 , \3319 , \3378 );
mand \mul_7_15/U$1117 ( \3380 , \3316 , \3379 );
mor \mul_7_15/U$1115 ( \3381 , \3315 , \3380 );
mand \mul_7_15/U$1112 ( \3382 , \3312 , \3381 );
mor \mul_7_15/U$1110 ( \3383 , \3311 , \3382 );
mand \mul_7_15/U$1107 ( \3384 , \3308 , \3383 );
mor \mul_7_15/U$1105 ( \3385 , \3307 , \3384 );
mand \mul_7_15/U$1102 ( \3386 , \3304 , \3385 );
mor \mul_7_15/U$1100 ( \3387 , \3303 , \3386 );
mand \mul_7_15/U$1097 ( \3388 , \3300 , \3387 );
mor \mul_7_15/U$1095 ( \3389 , \3299 , \3388 );
mand \mul_7_15/U$1092 ( \3390 , \3296 , \3389 );
mor \mul_7_15/U$1090 ( \3391 , \3295 , \3390 );
mand \mul_7_15/U$1073 ( \3392 , \2923_A[16] , \2997_B[5] );
mand \mul_7_15/U$994 ( \3393 , \3391 , \3392 );
mxor \mul_7_15/U$995 ( \3394 , \3391 , \3392 );
mxor \mul_7_15/U$1091 ( \3395 , \3296 , \3389 );
mand \mul_7_15/U$1074 ( \3396 , \2927_A[15] , \2997_B[5] );
mand \mul_7_15/U$999 ( \3397 , \3395 , \3396 );
mxor \mul_7_15/U$1000 ( \3398 , \3395 , \3396 );
mxor \mul_7_15/U$1096 ( \3399 , \3300 , \3387 );
mand \mul_7_15/U$1075 ( \3400 , \2931_A[14] , \2997_B[5] );
mand \mul_7_15/U$1004 ( \3401 , \3399 , \3400 );
mxor \mul_7_15/U$1005 ( \3402 , \3399 , \3400 );
mxor \mul_7_15/U$1101 ( \3403 , \3304 , \3385 );
mand \mul_7_15/U$1076 ( \3404 , \2935_A[13] , \2997_B[5] );
mand \mul_7_15/U$1009 ( \3405 , \3403 , \3404 );
mxor \mul_7_15/U$1010 ( \3406 , \3403 , \3404 );
mxor \mul_7_15/U$1106 ( \3407 , \3308 , \3383 );
mand \mul_7_15/U$1077 ( \3408 , \2939_A[12] , \2997_B[5] );
mand \mul_7_15/U$1014 ( \3409 , \3407 , \3408 );
mxor \mul_7_15/U$1015 ( \3410 , \3407 , \3408 );
mxor \mul_7_15/U$1111 ( \3411 , \3312 , \3381 );
mand \mul_7_15/U$1078 ( \3412 , \2943_A[11] , \2997_B[5] );
mand \mul_7_15/U$1019 ( \3413 , \3411 , \3412 );
mxor \mul_7_15/U$1020 ( \3414 , \3411 , \3412 );
mxor \mul_7_15/U$1116 ( \3415 , \3316 , \3379 );
mand \mul_7_15/U$1079 ( \3416 , \2947_A[10] , \2997_B[5] );
mand \mul_7_15/U$1024 ( \3417 , \3415 , \3416 );
mxor \mul_7_15/U$1025 ( \3418 , \3415 , \3416 );
mxor \mul_7_15/U$1121 ( \3419 , \3320 , \3377 );
mand \mul_7_15/U$1080 ( \3420 , \2951_A[9] , \2997_B[5] );
mand \mul_7_15/U$1029 ( \3421 , \3419 , \3420 );
mxor \mul_7_15/U$1030 ( \3422 , \3419 , \3420 );
mxor \mul_7_15/U$1126 ( \3423 , \3324 , \3375 );
mand \mul_7_15/U$1081 ( \3424 , \2955_A[8] , \2997_B[5] );
mand \mul_7_15/U$1034 ( \3425 , \3423 , \3424 );
mxor \mul_7_15/U$1035 ( \3426 , \3423 , \3424 );
mxor \mul_7_15/U$1131 ( \3427 , \3328 , \3373 );
mand \mul_7_15/U$1082 ( \3428 , \2959_A[7] , \2997_B[5] );
mand \mul_7_15/U$1039 ( \3429 , \3427 , \3428 );
mxor \mul_7_15/U$1040 ( \3430 , \3427 , \3428 );
mxor \mul_7_15/U$1136 ( \3431 , \3332 , \3371 );
mand \mul_7_15/U$1083 ( \3432 , \2963_A[6] , \2997_B[5] );
mand \mul_7_15/U$1044 ( \3433 , \3431 , \3432 );
mxor \mul_7_15/U$1045 ( \3434 , \3431 , \3432 );
mxor \mul_7_15/U$1141 ( \3435 , \3336 , \3369 );
mand \mul_7_15/U$1084 ( \3436 , \2967_A[5] , \2997_B[5] );
mand \mul_7_15/U$1049 ( \3437 , \3435 , \3436 );
mxor \mul_7_15/U$1050 ( \3438 , \3435 , \3436 );
mxor \mul_7_15/U$1146 ( \3439 , \3340 , \3367 );
mand \mul_7_15/U$1085 ( \3440 , \2971_A[4] , \2997_B[5] );
mand \mul_7_15/U$1054 ( \3441 , \3439 , \3440 );
mxor \mul_7_15/U$1055 ( \3442 , \3439 , \3440 );
mxor \mul_7_15/U$1151 ( \3443 , \3344 , \3365 );
mand \mul_7_15/U$1086 ( \3444 , \2975_A[3] , \2997_B[5] );
mand \mul_7_15/U$1059 ( \3445 , \3443 , \3444 );
mxor \mul_7_15/U$1060 ( \3446 , \3443 , \3444 );
mxor \mul_7_15/U$1156 ( \3447 , \3348 , \3363 );
mand \mul_7_15/U$1087 ( \3448 , \2979_A[2] , \2997_B[5] );
mand \mul_7_15/U$1064 ( \3449 , \3447 , \3448 );
mxor \mul_7_15/U$1065 ( \3450 , \3447 , \3448 );
mxor \mul_7_15/U$1161 ( \3451 , \3352 , \3361 );
mand \mul_7_15/U$1088 ( \3452 , \2983_A[1] , \2997_B[5] );
mand \mul_7_15/U$1069 ( \3453 , \3451 , \3452 );
mxor \mul_7_15/U$1070 ( \3454 , \3451 , \3452 );
mxor \mul_7_15/U$1166 ( \3455 , \3356 , \3359 );
mand \mul_7_15/U$1089 ( \3456 , \2986_A[0] , \2997_B[5] );
mand \mul_7_15/U$1071 ( \3457 , \3455 , \3456 );
mand \mul_7_15/U$1068 ( \3458 , \3454 , \3457 );
mor \mul_7_15/U$1066 ( \3459 , \3453 , \3458 );
mand \mul_7_15/U$1063 ( \3460 , \3450 , \3459 );
mor \mul_7_15/U$1061 ( \3461 , \3449 , \3460 );
mand \mul_7_15/U$1058 ( \3462 , \3446 , \3461 );
mor \mul_7_15/U$1056 ( \3463 , \3445 , \3462 );
mand \mul_7_15/U$1053 ( \3464 , \3442 , \3463 );
mor \mul_7_15/U$1051 ( \3465 , \3441 , \3464 );
mand \mul_7_15/U$1048 ( \3466 , \3438 , \3465 );
mor \mul_7_15/U$1046 ( \3467 , \3437 , \3466 );
mand \mul_7_15/U$1043 ( \3468 , \3434 , \3467 );
mor \mul_7_15/U$1041 ( \3469 , \3433 , \3468 );
mand \mul_7_15/U$1038 ( \3470 , \3430 , \3469 );
mor \mul_7_15/U$1036 ( \3471 , \3429 , \3470 );
mand \mul_7_15/U$1033 ( \3472 , \3426 , \3471 );
mor \mul_7_15/U$1031 ( \3473 , \3425 , \3472 );
mand \mul_7_15/U$1028 ( \3474 , \3422 , \3473 );
mor \mul_7_15/U$1026 ( \3475 , \3421 , \3474 );
mand \mul_7_15/U$1023 ( \3476 , \3418 , \3475 );
mor \mul_7_15/U$1021 ( \3477 , \3417 , \3476 );
mand \mul_7_15/U$1018 ( \3478 , \3414 , \3477 );
mor \mul_7_15/U$1016 ( \3479 , \3413 , \3478 );
mand \mul_7_15/U$1013 ( \3480 , \3410 , \3479 );
mor \mul_7_15/U$1011 ( \3481 , \3409 , \3480 );
mand \mul_7_15/U$1008 ( \3482 , \3406 , \3481 );
mor \mul_7_15/U$1006 ( \3483 , \3405 , \3482 );
mand \mul_7_15/U$1003 ( \3484 , \3402 , \3483 );
mor \mul_7_15/U$1001 ( \3485 , \3401 , \3484 );
mand \mul_7_15/U$998 ( \3486 , \3398 , \3485 );
mor \mul_7_15/U$996 ( \3487 , \3397 , \3486 );
mand \mul_7_15/U$993 ( \3488 , \3394 , \3487 );
mor \mul_7_15/U$991 ( \3489 , \3393 , \3488 );
mand \mul_7_15/U$974 ( \3490 , \2923_A[16] , \2996_B[6] );
mand \mul_7_15/U$895 ( \3491 , \3489 , \3490 );
mxor \mul_7_15/U$896 ( \3492 , \3489 , \3490 );
mxor \mul_7_15/U$992 ( \3493 , \3394 , \3487 );
mand \mul_7_15/U$975 ( \3494 , \2927_A[15] , \2996_B[6] );
mand \mul_7_15/U$900 ( \3495 , \3493 , \3494 );
mxor \mul_7_15/U$901 ( \3496 , \3493 , \3494 );
mxor \mul_7_15/U$997 ( \3497 , \3398 , \3485 );
mand \mul_7_15/U$976 ( \3498 , \2931_A[14] , \2996_B[6] );
mand \mul_7_15/U$905 ( \3499 , \3497 , \3498 );
mxor \mul_7_15/U$906 ( \3500 , \3497 , \3498 );
mxor \mul_7_15/U$1002 ( \3501 , \3402 , \3483 );
mand \mul_7_15/U$977 ( \3502 , \2935_A[13] , \2996_B[6] );
mand \mul_7_15/U$910 ( \3503 , \3501 , \3502 );
mxor \mul_7_15/U$911 ( \3504 , \3501 , \3502 );
mxor \mul_7_15/U$1007 ( \3505 , \3406 , \3481 );
mand \mul_7_15/U$978 ( \3506 , \2939_A[12] , \2996_B[6] );
mand \mul_7_15/U$915 ( \3507 , \3505 , \3506 );
mxor \mul_7_15/U$916 ( \3508 , \3505 , \3506 );
mxor \mul_7_15/U$1012 ( \3509 , \3410 , \3479 );
mand \mul_7_15/U$979 ( \3510 , \2943_A[11] , \2996_B[6] );
mand \mul_7_15/U$920 ( \3511 , \3509 , \3510 );
mxor \mul_7_15/U$921 ( \3512 , \3509 , \3510 );
mxor \mul_7_15/U$1017 ( \3513 , \3414 , \3477 );
mand \mul_7_15/U$980 ( \3514 , \2947_A[10] , \2996_B[6] );
mand \mul_7_15/U$925 ( \3515 , \3513 , \3514 );
mxor \mul_7_15/U$926 ( \3516 , \3513 , \3514 );
mxor \mul_7_15/U$1022 ( \3517 , \3418 , \3475 );
mand \mul_7_15/U$981 ( \3518 , \2951_A[9] , \2996_B[6] );
mand \mul_7_15/U$930 ( \3519 , \3517 , \3518 );
mxor \mul_7_15/U$931 ( \3520 , \3517 , \3518 );
mxor \mul_7_15/U$1027 ( \3521 , \3422 , \3473 );
mand \mul_7_15/U$982 ( \3522 , \2955_A[8] , \2996_B[6] );
mand \mul_7_15/U$935 ( \3523 , \3521 , \3522 );
mxor \mul_7_15/U$936 ( \3524 , \3521 , \3522 );
mxor \mul_7_15/U$1032 ( \3525 , \3426 , \3471 );
mand \mul_7_15/U$983 ( \3526 , \2959_A[7] , \2996_B[6] );
mand \mul_7_15/U$940 ( \3527 , \3525 , \3526 );
mxor \mul_7_15/U$941 ( \3528 , \3525 , \3526 );
mxor \mul_7_15/U$1037 ( \3529 , \3430 , \3469 );
mand \mul_7_15/U$984 ( \3530 , \2963_A[6] , \2996_B[6] );
mand \mul_7_15/U$945 ( \3531 , \3529 , \3530 );
mxor \mul_7_15/U$946 ( \3532 , \3529 , \3530 );
mxor \mul_7_15/U$1042 ( \3533 , \3434 , \3467 );
mand \mul_7_15/U$985 ( \3534 , \2967_A[5] , \2996_B[6] );
mand \mul_7_15/U$950 ( \3535 , \3533 , \3534 );
mxor \mul_7_15/U$951 ( \3536 , \3533 , \3534 );
mxor \mul_7_15/U$1047 ( \3537 , \3438 , \3465 );
mand \mul_7_15/U$986 ( \3538 , \2971_A[4] , \2996_B[6] );
mand \mul_7_15/U$955 ( \3539 , \3537 , \3538 );
mxor \mul_7_15/U$956 ( \3540 , \3537 , \3538 );
mxor \mul_7_15/U$1052 ( \3541 , \3442 , \3463 );
mand \mul_7_15/U$987 ( \3542 , \2975_A[3] , \2996_B[6] );
mand \mul_7_15/U$960 ( \3543 , \3541 , \3542 );
mxor \mul_7_15/U$961 ( \3544 , \3541 , \3542 );
mxor \mul_7_15/U$1057 ( \3545 , \3446 , \3461 );
mand \mul_7_15/U$988 ( \3546 , \2979_A[2] , \2996_B[6] );
mand \mul_7_15/U$965 ( \3547 , \3545 , \3546 );
mxor \mul_7_15/U$966 ( \3548 , \3545 , \3546 );
mxor \mul_7_15/U$1062 ( \3549 , \3450 , \3459 );
mand \mul_7_15/U$989 ( \3550 , \2983_A[1] , \2996_B[6] );
mand \mul_7_15/U$970 ( \3551 , \3549 , \3550 );
mxor \mul_7_15/U$971 ( \3552 , \3549 , \3550 );
mxor \mul_7_15/U$1067 ( \3553 , \3454 , \3457 );
mand \mul_7_15/U$990 ( \3554 , \2986_A[0] , \2996_B[6] );
mand \mul_7_15/U$972 ( \3555 , \3553 , \3554 );
mand \mul_7_15/U$969 ( \3556 , \3552 , \3555 );
mor \mul_7_15/U$967 ( \3557 , \3551 , \3556 );
mand \mul_7_15/U$964 ( \3558 , \3548 , \3557 );
mor \mul_7_15/U$962 ( \3559 , \3547 , \3558 );
mand \mul_7_15/U$959 ( \3560 , \3544 , \3559 );
mor \mul_7_15/U$957 ( \3561 , \3543 , \3560 );
mand \mul_7_15/U$954 ( \3562 , \3540 , \3561 );
mor \mul_7_15/U$952 ( \3563 , \3539 , \3562 );
mand \mul_7_15/U$949 ( \3564 , \3536 , \3563 );
mor \mul_7_15/U$947 ( \3565 , \3535 , \3564 );
mand \mul_7_15/U$944 ( \3566 , \3532 , \3565 );
mor \mul_7_15/U$942 ( \3567 , \3531 , \3566 );
mand \mul_7_15/U$939 ( \3568 , \3528 , \3567 );
mor \mul_7_15/U$937 ( \3569 , \3527 , \3568 );
mand \mul_7_15/U$934 ( \3570 , \3524 , \3569 );
mor \mul_7_15/U$932 ( \3571 , \3523 , \3570 );
mand \mul_7_15/U$929 ( \3572 , \3520 , \3571 );
mor \mul_7_15/U$927 ( \3573 , \3519 , \3572 );
mand \mul_7_15/U$924 ( \3574 , \3516 , \3573 );
mor \mul_7_15/U$922 ( \3575 , \3515 , \3574 );
mand \mul_7_15/U$919 ( \3576 , \3512 , \3575 );
mor \mul_7_15/U$917 ( \3577 , \3511 , \3576 );
mand \mul_7_15/U$914 ( \3578 , \3508 , \3577 );
mor \mul_7_15/U$912 ( \3579 , \3507 , \3578 );
mand \mul_7_15/U$909 ( \3580 , \3504 , \3579 );
mor \mul_7_15/U$907 ( \3581 , \3503 , \3580 );
mand \mul_7_15/U$904 ( \3582 , \3500 , \3581 );
mor \mul_7_15/U$902 ( \3583 , \3499 , \3582 );
mand \mul_7_15/U$899 ( \3584 , \3496 , \3583 );
mor \mul_7_15/U$897 ( \3585 , \3495 , \3584 );
mand \mul_7_15/U$894 ( \3586 , \3492 , \3585 );
mor \mul_7_15/U$892 ( \3587 , \3491 , \3586 );
mand \mul_7_15/U$875 ( \3588 , \2923_A[16] , \2995_B[7] );
mand \mul_7_15/U$796 ( \3589 , \3587 , \3588 );
mxor \mul_7_15/U$797 ( \3590 , \3587 , \3588 );
mxor \mul_7_15/U$893 ( \3591 , \3492 , \3585 );
mand \mul_7_15/U$876 ( \3592 , \2927_A[15] , \2995_B[7] );
mand \mul_7_15/U$801 ( \3593 , \3591 , \3592 );
mxor \mul_7_15/U$802 ( \3594 , \3591 , \3592 );
mxor \mul_7_15/U$898 ( \3595 , \3496 , \3583 );
mand \mul_7_15/U$877 ( \3596 , \2931_A[14] , \2995_B[7] );
mand \mul_7_15/U$806 ( \3597 , \3595 , \3596 );
mxor \mul_7_15/U$807 ( \3598 , \3595 , \3596 );
mxor \mul_7_15/U$903 ( \3599 , \3500 , \3581 );
mand \mul_7_15/U$878 ( \3600 , \2935_A[13] , \2995_B[7] );
mand \mul_7_15/U$811 ( \3601 , \3599 , \3600 );
mxor \mul_7_15/U$812 ( \3602 , \3599 , \3600 );
mxor \mul_7_15/U$908 ( \3603 , \3504 , \3579 );
mand \mul_7_15/U$879 ( \3604 , \2939_A[12] , \2995_B[7] );
mand \mul_7_15/U$816 ( \3605 , \3603 , \3604 );
mxor \mul_7_15/U$817 ( \3606 , \3603 , \3604 );
mxor \mul_7_15/U$913 ( \3607 , \3508 , \3577 );
mand \mul_7_15/U$880 ( \3608 , \2943_A[11] , \2995_B[7] );
mand \mul_7_15/U$821 ( \3609 , \3607 , \3608 );
mxor \mul_7_15/U$822 ( \3610 , \3607 , \3608 );
mxor \mul_7_15/U$918 ( \3611 , \3512 , \3575 );
mand \mul_7_15/U$881 ( \3612 , \2947_A[10] , \2995_B[7] );
mand \mul_7_15/U$826 ( \3613 , \3611 , \3612 );
mxor \mul_7_15/U$827 ( \3614 , \3611 , \3612 );
mxor \mul_7_15/U$923 ( \3615 , \3516 , \3573 );
mand \mul_7_15/U$882 ( \3616 , \2951_A[9] , \2995_B[7] );
mand \mul_7_15/U$831 ( \3617 , \3615 , \3616 );
mxor \mul_7_15/U$832 ( \3618 , \3615 , \3616 );
mxor \mul_7_15/U$928 ( \3619 , \3520 , \3571 );
mand \mul_7_15/U$883 ( \3620 , \2955_A[8] , \2995_B[7] );
mand \mul_7_15/U$836 ( \3621 , \3619 , \3620 );
mxor \mul_7_15/U$837 ( \3622 , \3619 , \3620 );
mxor \mul_7_15/U$933 ( \3623 , \3524 , \3569 );
mand \mul_7_15/U$884 ( \3624 , \2959_A[7] , \2995_B[7] );
mand \mul_7_15/U$841 ( \3625 , \3623 , \3624 );
mxor \mul_7_15/U$842 ( \3626 , \3623 , \3624 );
mxor \mul_7_15/U$938 ( \3627 , \3528 , \3567 );
mand \mul_7_15/U$885 ( \3628 , \2963_A[6] , \2995_B[7] );
mand \mul_7_15/U$846 ( \3629 , \3627 , \3628 );
mxor \mul_7_15/U$847 ( \3630 , \3627 , \3628 );
mxor \mul_7_15/U$943 ( \3631 , \3532 , \3565 );
mand \mul_7_15/U$886 ( \3632 , \2967_A[5] , \2995_B[7] );
mand \mul_7_15/U$851 ( \3633 , \3631 , \3632 );
mxor \mul_7_15/U$852 ( \3634 , \3631 , \3632 );
mxor \mul_7_15/U$948 ( \3635 , \3536 , \3563 );
mand \mul_7_15/U$887 ( \3636 , \2971_A[4] , \2995_B[7] );
mand \mul_7_15/U$856 ( \3637 , \3635 , \3636 );
mxor \mul_7_15/U$857 ( \3638 , \3635 , \3636 );
mxor \mul_7_15/U$953 ( \3639 , \3540 , \3561 );
mand \mul_7_15/U$888 ( \3640 , \2975_A[3] , \2995_B[7] );
mand \mul_7_15/U$861 ( \3641 , \3639 , \3640 );
mxor \mul_7_15/U$862 ( \3642 , \3639 , \3640 );
mxor \mul_7_15/U$958 ( \3643 , \3544 , \3559 );
mand \mul_7_15/U$889 ( \3644 , \2979_A[2] , \2995_B[7] );
mand \mul_7_15/U$866 ( \3645 , \3643 , \3644 );
mxor \mul_7_15/U$867 ( \3646 , \3643 , \3644 );
mxor \mul_7_15/U$963 ( \3647 , \3548 , \3557 );
mand \mul_7_15/U$890 ( \3648 , \2983_A[1] , \2995_B[7] );
mand \mul_7_15/U$871 ( \3649 , \3647 , \3648 );
mxor \mul_7_15/U$872 ( \3650 , \3647 , \3648 );
mxor \mul_7_15/U$968 ( \3651 , \3552 , \3555 );
mand \mul_7_15/U$891 ( \3652 , \2986_A[0] , \2995_B[7] );
mand \mul_7_15/U$873 ( \3653 , \3651 , \3652 );
mand \mul_7_15/U$870 ( \3654 , \3650 , \3653 );
mor \mul_7_15/U$868 ( \3655 , \3649 , \3654 );
mand \mul_7_15/U$865 ( \3656 , \3646 , \3655 );
mor \mul_7_15/U$863 ( \3657 , \3645 , \3656 );
mand \mul_7_15/U$860 ( \3658 , \3642 , \3657 );
mor \mul_7_15/U$858 ( \3659 , \3641 , \3658 );
mand \mul_7_15/U$855 ( \3660 , \3638 , \3659 );
mor \mul_7_15/U$853 ( \3661 , \3637 , \3660 );
mand \mul_7_15/U$850 ( \3662 , \3634 , \3661 );
mor \mul_7_15/U$848 ( \3663 , \3633 , \3662 );
mand \mul_7_15/U$845 ( \3664 , \3630 , \3663 );
mor \mul_7_15/U$843 ( \3665 , \3629 , \3664 );
mand \mul_7_15/U$840 ( \3666 , \3626 , \3665 );
mor \mul_7_15/U$838 ( \3667 , \3625 , \3666 );
mand \mul_7_15/U$835 ( \3668 , \3622 , \3667 );
mor \mul_7_15/U$833 ( \3669 , \3621 , \3668 );
mand \mul_7_15/U$830 ( \3670 , \3618 , \3669 );
mor \mul_7_15/U$828 ( \3671 , \3617 , \3670 );
mand \mul_7_15/U$825 ( \3672 , \3614 , \3671 );
mor \mul_7_15/U$823 ( \3673 , \3613 , \3672 );
mand \mul_7_15/U$820 ( \3674 , \3610 , \3673 );
mor \mul_7_15/U$818 ( \3675 , \3609 , \3674 );
mand \mul_7_15/U$815 ( \3676 , \3606 , \3675 );
mor \mul_7_15/U$813 ( \3677 , \3605 , \3676 );
mand \mul_7_15/U$810 ( \3678 , \3602 , \3677 );
mor \mul_7_15/U$808 ( \3679 , \3601 , \3678 );
mand \mul_7_15/U$805 ( \3680 , \3598 , \3679 );
mor \mul_7_15/U$803 ( \3681 , \3597 , \3680 );
mand \mul_7_15/U$800 ( \3682 , \3594 , \3681 );
mor \mul_7_15/U$798 ( \3683 , \3593 , \3682 );
mand \mul_7_15/U$795 ( \3684 , \3590 , \3683 );
mor \mul_7_15/U$793 ( \3685 , \3589 , \3684 );
mand \mul_7_15/U$776 ( \3686 , \2923_A[16] , \2994_B[8] );
mand \mul_7_15/U$697 ( \3687 , \3685 , \3686 );
mxor \mul_7_15/U$698 ( \3688 , \3685 , \3686 );
mxor \mul_7_15/U$794 ( \3689 , \3590 , \3683 );
mand \mul_7_15/U$777 ( \3690 , \2927_A[15] , \2994_B[8] );
mand \mul_7_15/U$702 ( \3691 , \3689 , \3690 );
mxor \mul_7_15/U$703 ( \3692 , \3689 , \3690 );
mxor \mul_7_15/U$799 ( \3693 , \3594 , \3681 );
mand \mul_7_15/U$778 ( \3694 , \2931_A[14] , \2994_B[8] );
mand \mul_7_15/U$707 ( \3695 , \3693 , \3694 );
mxor \mul_7_15/U$708 ( \3696 , \3693 , \3694 );
mxor \mul_7_15/U$804 ( \3697 , \3598 , \3679 );
mand \mul_7_15/U$779 ( \3698 , \2935_A[13] , \2994_B[8] );
mand \mul_7_15/U$712 ( \3699 , \3697 , \3698 );
mxor \mul_7_15/U$713 ( \3700 , \3697 , \3698 );
mxor \mul_7_15/U$809 ( \3701 , \3602 , \3677 );
mand \mul_7_15/U$780 ( \3702 , \2939_A[12] , \2994_B[8] );
mand \mul_7_15/U$717 ( \3703 , \3701 , \3702 );
mxor \mul_7_15/U$718 ( \3704 , \3701 , \3702 );
mxor \mul_7_15/U$814 ( \3705 , \3606 , \3675 );
mand \mul_7_15/U$781 ( \3706 , \2943_A[11] , \2994_B[8] );
mand \mul_7_15/U$722 ( \3707 , \3705 , \3706 );
mxor \mul_7_15/U$723 ( \3708 , \3705 , \3706 );
mxor \mul_7_15/U$819 ( \3709 , \3610 , \3673 );
mand \mul_7_15/U$782 ( \3710 , \2947_A[10] , \2994_B[8] );
mand \mul_7_15/U$727 ( \3711 , \3709 , \3710 );
mxor \mul_7_15/U$728 ( \3712 , \3709 , \3710 );
mxor \mul_7_15/U$824 ( \3713 , \3614 , \3671 );
mand \mul_7_15/U$783 ( \3714 , \2951_A[9] , \2994_B[8] );
mand \mul_7_15/U$732 ( \3715 , \3713 , \3714 );
mxor \mul_7_15/U$733 ( \3716 , \3713 , \3714 );
mxor \mul_7_15/U$829 ( \3717 , \3618 , \3669 );
mand \mul_7_15/U$784 ( \3718 , \2955_A[8] , \2994_B[8] );
mand \mul_7_15/U$737 ( \3719 , \3717 , \3718 );
mxor \mul_7_15/U$738 ( \3720 , \3717 , \3718 );
mxor \mul_7_15/U$834 ( \3721 , \3622 , \3667 );
mand \mul_7_15/U$785 ( \3722 , \2959_A[7] , \2994_B[8] );
mand \mul_7_15/U$742 ( \3723 , \3721 , \3722 );
mxor \mul_7_15/U$743 ( \3724 , \3721 , \3722 );
mxor \mul_7_15/U$839 ( \3725 , \3626 , \3665 );
mand \mul_7_15/U$786 ( \3726 , \2963_A[6] , \2994_B[8] );
mand \mul_7_15/U$747 ( \3727 , \3725 , \3726 );
mxor \mul_7_15/U$748 ( \3728 , \3725 , \3726 );
mxor \mul_7_15/U$844 ( \3729 , \3630 , \3663 );
mand \mul_7_15/U$787 ( \3730 , \2967_A[5] , \2994_B[8] );
mand \mul_7_15/U$752 ( \3731 , \3729 , \3730 );
mxor \mul_7_15/U$753 ( \3732 , \3729 , \3730 );
mxor \mul_7_15/U$849 ( \3733 , \3634 , \3661 );
mand \mul_7_15/U$788 ( \3734 , \2971_A[4] , \2994_B[8] );
mand \mul_7_15/U$757 ( \3735 , \3733 , \3734 );
mxor \mul_7_15/U$758 ( \3736 , \3733 , \3734 );
mxor \mul_7_15/U$854 ( \3737 , \3638 , \3659 );
mand \mul_7_15/U$789 ( \3738 , \2975_A[3] , \2994_B[8] );
mand \mul_7_15/U$762 ( \3739 , \3737 , \3738 );
mxor \mul_7_15/U$763 ( \3740 , \3737 , \3738 );
mxor \mul_7_15/U$859 ( \3741 , \3642 , \3657 );
mand \mul_7_15/U$790 ( \3742 , \2979_A[2] , \2994_B[8] );
mand \mul_7_15/U$767 ( \3743 , \3741 , \3742 );
mxor \mul_7_15/U$768 ( \3744 , \3741 , \3742 );
mxor \mul_7_15/U$864 ( \3745 , \3646 , \3655 );
mand \mul_7_15/U$791 ( \3746 , \2983_A[1] , \2994_B[8] );
mand \mul_7_15/U$772 ( \3747 , \3745 , \3746 );
mxor \mul_7_15/U$773 ( \3748 , \3745 , \3746 );
mxor \mul_7_15/U$869 ( \3749 , \3650 , \3653 );
mand \mul_7_15/U$792 ( \3750 , \2986_A[0] , \2994_B[8] );
mand \mul_7_15/U$774 ( \3751 , \3749 , \3750 );
mand \mul_7_15/U$771 ( \3752 , \3748 , \3751 );
mor \mul_7_15/U$769 ( \3753 , \3747 , \3752 );
mand \mul_7_15/U$766 ( \3754 , \3744 , \3753 );
mor \mul_7_15/U$764 ( \3755 , \3743 , \3754 );
mand \mul_7_15/U$761 ( \3756 , \3740 , \3755 );
mor \mul_7_15/U$759 ( \3757 , \3739 , \3756 );
mand \mul_7_15/U$756 ( \3758 , \3736 , \3757 );
mor \mul_7_15/U$754 ( \3759 , \3735 , \3758 );
mand \mul_7_15/U$751 ( \3760 , \3732 , \3759 );
mor \mul_7_15/U$749 ( \3761 , \3731 , \3760 );
mand \mul_7_15/U$746 ( \3762 , \3728 , \3761 );
mor \mul_7_15/U$744 ( \3763 , \3727 , \3762 );
mand \mul_7_15/U$741 ( \3764 , \3724 , \3763 );
mor \mul_7_15/U$739 ( \3765 , \3723 , \3764 );
mand \mul_7_15/U$736 ( \3766 , \3720 , \3765 );
mor \mul_7_15/U$734 ( \3767 , \3719 , \3766 );
mand \mul_7_15/U$731 ( \3768 , \3716 , \3767 );
mor \mul_7_15/U$729 ( \3769 , \3715 , \3768 );
mand \mul_7_15/U$726 ( \3770 , \3712 , \3769 );
mor \mul_7_15/U$724 ( \3771 , \3711 , \3770 );
mand \mul_7_15/U$721 ( \3772 , \3708 , \3771 );
mor \mul_7_15/U$719 ( \3773 , \3707 , \3772 );
mand \mul_7_15/U$716 ( \3774 , \3704 , \3773 );
mor \mul_7_15/U$714 ( \3775 , \3703 , \3774 );
mand \mul_7_15/U$711 ( \3776 , \3700 , \3775 );
mor \mul_7_15/U$709 ( \3777 , \3699 , \3776 );
mand \mul_7_15/U$706 ( \3778 , \3696 , \3777 );
mor \mul_7_15/U$704 ( \3779 , \3695 , \3778 );
mand \mul_7_15/U$701 ( \3780 , \3692 , \3779 );
mor \mul_7_15/U$699 ( \3781 , \3691 , \3780 );
mand \mul_7_15/U$696 ( \3782 , \3688 , \3781 );
mor \mul_7_15/U$694 ( \3783 , \3687 , \3782 );
mand \mul_7_15/U$677 ( \3784 , \2923_A[16] , \2993_B[9] );
mand \mul_7_15/U$598 ( \3785 , \3783 , \3784 );
mxor \mul_7_15/U$599 ( \3786 , \3783 , \3784 );
mxor \mul_7_15/U$695 ( \3787 , \3688 , \3781 );
mand \mul_7_15/U$678 ( \3788 , \2927_A[15] , \2993_B[9] );
mand \mul_7_15/U$603 ( \3789 , \3787 , \3788 );
mxor \mul_7_15/U$604 ( \3790 , \3787 , \3788 );
mxor \mul_7_15/U$700 ( \3791 , \3692 , \3779 );
mand \mul_7_15/U$679 ( \3792 , \2931_A[14] , \2993_B[9] );
mand \mul_7_15/U$608 ( \3793 , \3791 , \3792 );
mxor \mul_7_15/U$609 ( \3794 , \3791 , \3792 );
mxor \mul_7_15/U$705 ( \3795 , \3696 , \3777 );
mand \mul_7_15/U$680 ( \3796 , \2935_A[13] , \2993_B[9] );
mand \mul_7_15/U$613 ( \3797 , \3795 , \3796 );
mxor \mul_7_15/U$614 ( \3798 , \3795 , \3796 );
mxor \mul_7_15/U$710 ( \3799 , \3700 , \3775 );
mand \mul_7_15/U$681 ( \3800 , \2939_A[12] , \2993_B[9] );
mand \mul_7_15/U$618 ( \3801 , \3799 , \3800 );
mxor \mul_7_15/U$619 ( \3802 , \3799 , \3800 );
mxor \mul_7_15/U$715 ( \3803 , \3704 , \3773 );
mand \mul_7_15/U$682 ( \3804 , \2943_A[11] , \2993_B[9] );
mand \mul_7_15/U$623 ( \3805 , \3803 , \3804 );
mxor \mul_7_15/U$624 ( \3806 , \3803 , \3804 );
mxor \mul_7_15/U$720 ( \3807 , \3708 , \3771 );
mand \mul_7_15/U$683 ( \3808 , \2947_A[10] , \2993_B[9] );
mand \mul_7_15/U$628 ( \3809 , \3807 , \3808 );
mxor \mul_7_15/U$629 ( \3810 , \3807 , \3808 );
mxor \mul_7_15/U$725 ( \3811 , \3712 , \3769 );
mand \mul_7_15/U$684 ( \3812 , \2951_A[9] , \2993_B[9] );
mand \mul_7_15/U$633 ( \3813 , \3811 , \3812 );
mxor \mul_7_15/U$634 ( \3814 , \3811 , \3812 );
mxor \mul_7_15/U$730 ( \3815 , \3716 , \3767 );
mand \mul_7_15/U$685 ( \3816 , \2955_A[8] , \2993_B[9] );
mand \mul_7_15/U$638 ( \3817 , \3815 , \3816 );
mxor \mul_7_15/U$639 ( \3818 , \3815 , \3816 );
mxor \mul_7_15/U$735 ( \3819 , \3720 , \3765 );
mand \mul_7_15/U$686 ( \3820 , \2959_A[7] , \2993_B[9] );
mand \mul_7_15/U$643 ( \3821 , \3819 , \3820 );
mxor \mul_7_15/U$644 ( \3822 , \3819 , \3820 );
mxor \mul_7_15/U$740 ( \3823 , \3724 , \3763 );
mand \mul_7_15/U$687 ( \3824 , \2963_A[6] , \2993_B[9] );
mand \mul_7_15/U$648 ( \3825 , \3823 , \3824 );
mxor \mul_7_15/U$649 ( \3826 , \3823 , \3824 );
mxor \mul_7_15/U$745 ( \3827 , \3728 , \3761 );
mand \mul_7_15/U$688 ( \3828 , \2967_A[5] , \2993_B[9] );
mand \mul_7_15/U$653 ( \3829 , \3827 , \3828 );
mxor \mul_7_15/U$654 ( \3830 , \3827 , \3828 );
mxor \mul_7_15/U$750 ( \3831 , \3732 , \3759 );
mand \mul_7_15/U$689 ( \3832 , \2971_A[4] , \2993_B[9] );
mand \mul_7_15/U$658 ( \3833 , \3831 , \3832 );
mxor \mul_7_15/U$659 ( \3834 , \3831 , \3832 );
mxor \mul_7_15/U$755 ( \3835 , \3736 , \3757 );
mand \mul_7_15/U$690 ( \3836 , \2975_A[3] , \2993_B[9] );
mand \mul_7_15/U$663 ( \3837 , \3835 , \3836 );
mxor \mul_7_15/U$664 ( \3838 , \3835 , \3836 );
mxor \mul_7_15/U$760 ( \3839 , \3740 , \3755 );
mand \mul_7_15/U$691 ( \3840 , \2979_A[2] , \2993_B[9] );
mand \mul_7_15/U$668 ( \3841 , \3839 , \3840 );
mxor \mul_7_15/U$669 ( \3842 , \3839 , \3840 );
mxor \mul_7_15/U$765 ( \3843 , \3744 , \3753 );
mand \mul_7_15/U$692 ( \3844 , \2983_A[1] , \2993_B[9] );
mand \mul_7_15/U$673 ( \3845 , \3843 , \3844 );
mxor \mul_7_15/U$674 ( \3846 , \3843 , \3844 );
mxor \mul_7_15/U$770 ( \3847 , \3748 , \3751 );
mand \mul_7_15/U$693 ( \3848 , \2986_A[0] , \2993_B[9] );
mand \mul_7_15/U$675 ( \3849 , \3847 , \3848 );
mand \mul_7_15/U$672 ( \3850 , \3846 , \3849 );
mor \mul_7_15/U$670 ( \3851 , \3845 , \3850 );
mand \mul_7_15/U$667 ( \3852 , \3842 , \3851 );
mor \mul_7_15/U$665 ( \3853 , \3841 , \3852 );
mand \mul_7_15/U$662 ( \3854 , \3838 , \3853 );
mor \mul_7_15/U$660 ( \3855 , \3837 , \3854 );
mand \mul_7_15/U$657 ( \3856 , \3834 , \3855 );
mor \mul_7_15/U$655 ( \3857 , \3833 , \3856 );
mand \mul_7_15/U$652 ( \3858 , \3830 , \3857 );
mor \mul_7_15/U$650 ( \3859 , \3829 , \3858 );
mand \mul_7_15/U$647 ( \3860 , \3826 , \3859 );
mor \mul_7_15/U$645 ( \3861 , \3825 , \3860 );
mand \mul_7_15/U$642 ( \3862 , \3822 , \3861 );
mor \mul_7_15/U$640 ( \3863 , \3821 , \3862 );
mand \mul_7_15/U$637 ( \3864 , \3818 , \3863 );
mor \mul_7_15/U$635 ( \3865 , \3817 , \3864 );
mand \mul_7_15/U$632 ( \3866 , \3814 , \3865 );
mor \mul_7_15/U$630 ( \3867 , \3813 , \3866 );
mand \mul_7_15/U$627 ( \3868 , \3810 , \3867 );
mor \mul_7_15/U$625 ( \3869 , \3809 , \3868 );
mand \mul_7_15/U$622 ( \3870 , \3806 , \3869 );
mor \mul_7_15/U$620 ( \3871 , \3805 , \3870 );
mand \mul_7_15/U$617 ( \3872 , \3802 , \3871 );
mor \mul_7_15/U$615 ( \3873 , \3801 , \3872 );
mand \mul_7_15/U$612 ( \3874 , \3798 , \3873 );
mor \mul_7_15/U$610 ( \3875 , \3797 , \3874 );
mand \mul_7_15/U$607 ( \3876 , \3794 , \3875 );
mor \mul_7_15/U$605 ( \3877 , \3793 , \3876 );
mand \mul_7_15/U$602 ( \3878 , \3790 , \3877 );
mor \mul_7_15/U$600 ( \3879 , \3789 , \3878 );
mand \mul_7_15/U$597 ( \3880 , \3786 , \3879 );
mor \mul_7_15/U$595 ( \3881 , \3785 , \3880 );
mand \mul_7_15/U$578 ( \3882 , \2923_A[16] , \2992_B[10] );
mand \mul_7_15/U$499 ( \3883 , \3881 , \3882 );
mxor \mul_7_15/U$500 ( \3884 , \3881 , \3882 );
mxor \mul_7_15/U$596 ( \3885 , \3786 , \3879 );
mand \mul_7_15/U$579 ( \3886 , \2927_A[15] , \2992_B[10] );
mand \mul_7_15/U$504 ( \3887 , \3885 , \3886 );
mxor \mul_7_15/U$505 ( \3888 , \3885 , \3886 );
mxor \mul_7_15/U$601 ( \3889 , \3790 , \3877 );
mand \mul_7_15/U$580 ( \3890 , \2931_A[14] , \2992_B[10] );
mand \mul_7_15/U$509 ( \3891 , \3889 , \3890 );
mxor \mul_7_15/U$510 ( \3892 , \3889 , \3890 );
mxor \mul_7_15/U$606 ( \3893 , \3794 , \3875 );
mand \mul_7_15/U$581 ( \3894 , \2935_A[13] , \2992_B[10] );
mand \mul_7_15/U$514 ( \3895 , \3893 , \3894 );
mxor \mul_7_15/U$515 ( \3896 , \3893 , \3894 );
mxor \mul_7_15/U$611 ( \3897 , \3798 , \3873 );
mand \mul_7_15/U$582 ( \3898 , \2939_A[12] , \2992_B[10] );
mand \mul_7_15/U$519 ( \3899 , \3897 , \3898 );
mxor \mul_7_15/U$520 ( \3900 , \3897 , \3898 );
mxor \mul_7_15/U$616 ( \3901 , \3802 , \3871 );
mand \mul_7_15/U$583 ( \3902 , \2943_A[11] , \2992_B[10] );
mand \mul_7_15/U$524 ( \3903 , \3901 , \3902 );
mxor \mul_7_15/U$525 ( \3904 , \3901 , \3902 );
mxor \mul_7_15/U$621 ( \3905 , \3806 , \3869 );
mand \mul_7_15/U$584 ( \3906 , \2947_A[10] , \2992_B[10] );
mand \mul_7_15/U$529 ( \3907 , \3905 , \3906 );
mxor \mul_7_15/U$530 ( \3908 , \3905 , \3906 );
mxor \mul_7_15/U$626 ( \3909 , \3810 , \3867 );
mand \mul_7_15/U$585 ( \3910 , \2951_A[9] , \2992_B[10] );
mand \mul_7_15/U$534 ( \3911 , \3909 , \3910 );
mxor \mul_7_15/U$535 ( \3912 , \3909 , \3910 );
mxor \mul_7_15/U$631 ( \3913 , \3814 , \3865 );
mand \mul_7_15/U$586 ( \3914 , \2955_A[8] , \2992_B[10] );
mand \mul_7_15/U$539 ( \3915 , \3913 , \3914 );
mxor \mul_7_15/U$540 ( \3916 , \3913 , \3914 );
mxor \mul_7_15/U$636 ( \3917 , \3818 , \3863 );
mand \mul_7_15/U$587 ( \3918 , \2959_A[7] , \2992_B[10] );
mand \mul_7_15/U$544 ( \3919 , \3917 , \3918 );
mxor \mul_7_15/U$545 ( \3920 , \3917 , \3918 );
mxor \mul_7_15/U$641 ( \3921 , \3822 , \3861 );
mand \mul_7_15/U$588 ( \3922 , \2963_A[6] , \2992_B[10] );
mand \mul_7_15/U$549 ( \3923 , \3921 , \3922 );
mxor \mul_7_15/U$550 ( \3924 , \3921 , \3922 );
mxor \mul_7_15/U$646 ( \3925 , \3826 , \3859 );
mand \mul_7_15/U$589 ( \3926 , \2967_A[5] , \2992_B[10] );
mand \mul_7_15/U$554 ( \3927 , \3925 , \3926 );
mxor \mul_7_15/U$555 ( \3928 , \3925 , \3926 );
mxor \mul_7_15/U$651 ( \3929 , \3830 , \3857 );
mand \mul_7_15/U$590 ( \3930 , \2971_A[4] , \2992_B[10] );
mand \mul_7_15/U$559 ( \3931 , \3929 , \3930 );
mxor \mul_7_15/U$560 ( \3932 , \3929 , \3930 );
mxor \mul_7_15/U$656 ( \3933 , \3834 , \3855 );
mand \mul_7_15/U$591 ( \3934 , \2975_A[3] , \2992_B[10] );
mand \mul_7_15/U$564 ( \3935 , \3933 , \3934 );
mxor \mul_7_15/U$565 ( \3936 , \3933 , \3934 );
mxor \mul_7_15/U$661 ( \3937 , \3838 , \3853 );
mand \mul_7_15/U$592 ( \3938 , \2979_A[2] , \2992_B[10] );
mand \mul_7_15/U$569 ( \3939 , \3937 , \3938 );
mxor \mul_7_15/U$570 ( \3940 , \3937 , \3938 );
mxor \mul_7_15/U$666 ( \3941 , \3842 , \3851 );
mand \mul_7_15/U$593 ( \3942 , \2983_A[1] , \2992_B[10] );
mand \mul_7_15/U$574 ( \3943 , \3941 , \3942 );
mxor \mul_7_15/U$575 ( \3944 , \3941 , \3942 );
mxor \mul_7_15/U$671 ( \3945 , \3846 , \3849 );
mand \mul_7_15/U$594 ( \3946 , \2986_A[0] , \2992_B[10] );
mand \mul_7_15/U$576 ( \3947 , \3945 , \3946 );
mand \mul_7_15/U$573 ( \3948 , \3944 , \3947 );
mor \mul_7_15/U$571 ( \3949 , \3943 , \3948 );
mand \mul_7_15/U$568 ( \3950 , \3940 , \3949 );
mor \mul_7_15/U$566 ( \3951 , \3939 , \3950 );
mand \mul_7_15/U$563 ( \3952 , \3936 , \3951 );
mor \mul_7_15/U$561 ( \3953 , \3935 , \3952 );
mand \mul_7_15/U$558 ( \3954 , \3932 , \3953 );
mor \mul_7_15/U$556 ( \3955 , \3931 , \3954 );
mand \mul_7_15/U$553 ( \3956 , \3928 , \3955 );
mor \mul_7_15/U$551 ( \3957 , \3927 , \3956 );
mand \mul_7_15/U$548 ( \3958 , \3924 , \3957 );
mor \mul_7_15/U$546 ( \3959 , \3923 , \3958 );
mand \mul_7_15/U$543 ( \3960 , \3920 , \3959 );
mor \mul_7_15/U$541 ( \3961 , \3919 , \3960 );
mand \mul_7_15/U$538 ( \3962 , \3916 , \3961 );
mor \mul_7_15/U$536 ( \3963 , \3915 , \3962 );
mand \mul_7_15/U$533 ( \3964 , \3912 , \3963 );
mor \mul_7_15/U$531 ( \3965 , \3911 , \3964 );
mand \mul_7_15/U$528 ( \3966 , \3908 , \3965 );
mor \mul_7_15/U$526 ( \3967 , \3907 , \3966 );
mand \mul_7_15/U$523 ( \3968 , \3904 , \3967 );
mor \mul_7_15/U$521 ( \3969 , \3903 , \3968 );
mand \mul_7_15/U$518 ( \3970 , \3900 , \3969 );
mor \mul_7_15/U$516 ( \3971 , \3899 , \3970 );
mand \mul_7_15/U$513 ( \3972 , \3896 , \3971 );
mor \mul_7_15/U$511 ( \3973 , \3895 , \3972 );
mand \mul_7_15/U$508 ( \3974 , \3892 , \3973 );
mor \mul_7_15/U$506 ( \3975 , \3891 , \3974 );
mand \mul_7_15/U$503 ( \3976 , \3888 , \3975 );
mor \mul_7_15/U$501 ( \3977 , \3887 , \3976 );
mand \mul_7_15/U$498 ( \3978 , \3884 , \3977 );
mor \mul_7_15/U$496 ( \3979 , \3883 , \3978 );
mand \mul_7_15/U$479 ( \3980 , \2923_A[16] , \2991_B[11] );
mand \mul_7_15/U$400 ( \3981 , \3979 , \3980 );
mxor \mul_7_15/U$401 ( \3982 , \3979 , \3980 );
mxor \mul_7_15/U$497 ( \3983 , \3884 , \3977 );
mand \mul_7_15/U$480 ( \3984 , \2927_A[15] , \2991_B[11] );
mand \mul_7_15/U$405 ( \3985 , \3983 , \3984 );
mxor \mul_7_15/U$406 ( \3986 , \3983 , \3984 );
mxor \mul_7_15/U$502 ( \3987 , \3888 , \3975 );
mand \mul_7_15/U$481 ( \3988 , \2931_A[14] , \2991_B[11] );
mand \mul_7_15/U$410 ( \3989 , \3987 , \3988 );
mxor \mul_7_15/U$411 ( \3990 , \3987 , \3988 );
mxor \mul_7_15/U$507 ( \3991 , \3892 , \3973 );
mand \mul_7_15/U$482 ( \3992 , \2935_A[13] , \2991_B[11] );
mand \mul_7_15/U$415 ( \3993 , \3991 , \3992 );
mxor \mul_7_15/U$416 ( \3994 , \3991 , \3992 );
mxor \mul_7_15/U$512 ( \3995 , \3896 , \3971 );
mand \mul_7_15/U$483 ( \3996 , \2939_A[12] , \2991_B[11] );
mand \mul_7_15/U$420 ( \3997 , \3995 , \3996 );
mxor \mul_7_15/U$421 ( \3998 , \3995 , \3996 );
mxor \mul_7_15/U$517 ( \3999 , \3900 , \3969 );
mand \mul_7_15/U$484 ( \4000 , \2943_A[11] , \2991_B[11] );
mand \mul_7_15/U$425 ( \4001 , \3999 , \4000 );
mxor \mul_7_15/U$426 ( \4002 , \3999 , \4000 );
mxor \mul_7_15/U$522 ( \4003 , \3904 , \3967 );
mand \mul_7_15/U$485 ( \4004 , \2947_A[10] , \2991_B[11] );
mand \mul_7_15/U$430 ( \4005 , \4003 , \4004 );
mxor \mul_7_15/U$431 ( \4006 , \4003 , \4004 );
mxor \mul_7_15/U$527 ( \4007 , \3908 , \3965 );
mand \mul_7_15/U$486 ( \4008 , \2951_A[9] , \2991_B[11] );
mand \mul_7_15/U$435 ( \4009 , \4007 , \4008 );
mxor \mul_7_15/U$436 ( \4010 , \4007 , \4008 );
mxor \mul_7_15/U$532 ( \4011 , \3912 , \3963 );
mand \mul_7_15/U$487 ( \4012 , \2955_A[8] , \2991_B[11] );
mand \mul_7_15/U$440 ( \4013 , \4011 , \4012 );
mxor \mul_7_15/U$441 ( \4014 , \4011 , \4012 );
mxor \mul_7_15/U$537 ( \4015 , \3916 , \3961 );
mand \mul_7_15/U$488 ( \4016 , \2959_A[7] , \2991_B[11] );
mand \mul_7_15/U$445 ( \4017 , \4015 , \4016 );
mxor \mul_7_15/U$446 ( \4018 , \4015 , \4016 );
mxor \mul_7_15/U$542 ( \4019 , \3920 , \3959 );
mand \mul_7_15/U$489 ( \4020 , \2963_A[6] , \2991_B[11] );
mand \mul_7_15/U$450 ( \4021 , \4019 , \4020 );
mxor \mul_7_15/U$451 ( \4022 , \4019 , \4020 );
mxor \mul_7_15/U$547 ( \4023 , \3924 , \3957 );
mand \mul_7_15/U$490 ( \4024 , \2967_A[5] , \2991_B[11] );
mand \mul_7_15/U$455 ( \4025 , \4023 , \4024 );
mxor \mul_7_15/U$456 ( \4026 , \4023 , \4024 );
mxor \mul_7_15/U$552 ( \4027 , \3928 , \3955 );
mand \mul_7_15/U$491 ( \4028 , \2971_A[4] , \2991_B[11] );
mand \mul_7_15/U$460 ( \4029 , \4027 , \4028 );
mxor \mul_7_15/U$461 ( \4030 , \4027 , \4028 );
mxor \mul_7_15/U$557 ( \4031 , \3932 , \3953 );
mand \mul_7_15/U$492 ( \4032 , \2975_A[3] , \2991_B[11] );
mand \mul_7_15/U$465 ( \4033 , \4031 , \4032 );
mxor \mul_7_15/U$466 ( \4034 , \4031 , \4032 );
mxor \mul_7_15/U$562 ( \4035 , \3936 , \3951 );
mand \mul_7_15/U$493 ( \4036 , \2979_A[2] , \2991_B[11] );
mand \mul_7_15/U$470 ( \4037 , \4035 , \4036 );
mxor \mul_7_15/U$471 ( \4038 , \4035 , \4036 );
mxor \mul_7_15/U$567 ( \4039 , \3940 , \3949 );
mand \mul_7_15/U$494 ( \4040 , \2983_A[1] , \2991_B[11] );
mand \mul_7_15/U$475 ( \4041 , \4039 , \4040 );
mxor \mul_7_15/U$476 ( \4042 , \4039 , \4040 );
mxor \mul_7_15/U$572 ( \4043 , \3944 , \3947 );
mand \mul_7_15/U$495 ( \4044 , \2986_A[0] , \2991_B[11] );
mand \mul_7_15/U$477 ( \4045 , \4043 , \4044 );
mand \mul_7_15/U$474 ( \4046 , \4042 , \4045 );
mor \mul_7_15/U$472 ( \4047 , \4041 , \4046 );
mand \mul_7_15/U$469 ( \4048 , \4038 , \4047 );
mor \mul_7_15/U$467 ( \4049 , \4037 , \4048 );
mand \mul_7_15/U$464 ( \4050 , \4034 , \4049 );
mor \mul_7_15/U$462 ( \4051 , \4033 , \4050 );
mand \mul_7_15/U$459 ( \4052 , \4030 , \4051 );
mor \mul_7_15/U$457 ( \4053 , \4029 , \4052 );
mand \mul_7_15/U$454 ( \4054 , \4026 , \4053 );
mor \mul_7_15/U$452 ( \4055 , \4025 , \4054 );
mand \mul_7_15/U$449 ( \4056 , \4022 , \4055 );
mor \mul_7_15/U$447 ( \4057 , \4021 , \4056 );
mand \mul_7_15/U$444 ( \4058 , \4018 , \4057 );
mor \mul_7_15/U$442 ( \4059 , \4017 , \4058 );
mand \mul_7_15/U$439 ( \4060 , \4014 , \4059 );
mor \mul_7_15/U$437 ( \4061 , \4013 , \4060 );
mand \mul_7_15/U$434 ( \4062 , \4010 , \4061 );
mor \mul_7_15/U$432 ( \4063 , \4009 , \4062 );
mand \mul_7_15/U$429 ( \4064 , \4006 , \4063 );
mor \mul_7_15/U$427 ( \4065 , \4005 , \4064 );
mand \mul_7_15/U$424 ( \4066 , \4002 , \4065 );
mor \mul_7_15/U$422 ( \4067 , \4001 , \4066 );
mand \mul_7_15/U$419 ( \4068 , \3998 , \4067 );
mor \mul_7_15/U$417 ( \4069 , \3997 , \4068 );
mand \mul_7_15/U$414 ( \4070 , \3994 , \4069 );
mor \mul_7_15/U$412 ( \4071 , \3993 , \4070 );
mand \mul_7_15/U$409 ( \4072 , \3990 , \4071 );
mor \mul_7_15/U$407 ( \4073 , \3989 , \4072 );
mand \mul_7_15/U$404 ( \4074 , \3986 , \4073 );
mor \mul_7_15/U$402 ( \4075 , \3985 , \4074 );
mand \mul_7_15/U$399 ( \4076 , \3982 , \4075 );
mor \mul_7_15/U$397 ( \4077 , \3981 , \4076 );
mand \mul_7_15/U$380 ( \4078 , \2923_A[16] , \2990_B[12] );
mand \mul_7_15/U$301 ( \4079 , \4077 , \4078 );
mxor \mul_7_15/U$302 ( \4080 , \4077 , \4078 );
mxor \mul_7_15/U$398 ( \4081 , \3982 , \4075 );
mand \mul_7_15/U$381 ( \4082 , \2927_A[15] , \2990_B[12] );
mand \mul_7_15/U$306 ( \4083 , \4081 , \4082 );
mxor \mul_7_15/U$307 ( \4084 , \4081 , \4082 );
mxor \mul_7_15/U$403 ( \4085 , \3986 , \4073 );
mand \mul_7_15/U$382 ( \4086 , \2931_A[14] , \2990_B[12] );
mand \mul_7_15/U$311 ( \4087 , \4085 , \4086 );
mxor \mul_7_15/U$312 ( \4088 , \4085 , \4086 );
mxor \mul_7_15/U$408 ( \4089 , \3990 , \4071 );
mand \mul_7_15/U$383 ( \4090 , \2935_A[13] , \2990_B[12] );
mand \mul_7_15/U$316 ( \4091 , \4089 , \4090 );
mxor \mul_7_15/U$317 ( \4092 , \4089 , \4090 );
mxor \mul_7_15/U$413 ( \4093 , \3994 , \4069 );
mand \mul_7_15/U$384 ( \4094 , \2939_A[12] , \2990_B[12] );
mand \mul_7_15/U$321 ( \4095 , \4093 , \4094 );
mxor \mul_7_15/U$322 ( \4096 , \4093 , \4094 );
mxor \mul_7_15/U$418 ( \4097 , \3998 , \4067 );
mand \mul_7_15/U$385 ( \4098 , \2943_A[11] , \2990_B[12] );
mand \mul_7_15/U$326 ( \4099 , \4097 , \4098 );
mxor \mul_7_15/U$327 ( \4100 , \4097 , \4098 );
mxor \mul_7_15/U$423 ( \4101 , \4002 , \4065 );
mand \mul_7_15/U$386 ( \4102 , \2947_A[10] , \2990_B[12] );
mand \mul_7_15/U$331 ( \4103 , \4101 , \4102 );
mxor \mul_7_15/U$332 ( \4104 , \4101 , \4102 );
mxor \mul_7_15/U$428 ( \4105 , \4006 , \4063 );
mand \mul_7_15/U$387 ( \4106 , \2951_A[9] , \2990_B[12] );
mand \mul_7_15/U$336 ( \4107 , \4105 , \4106 );
mxor \mul_7_15/U$337 ( \4108 , \4105 , \4106 );
mxor \mul_7_15/U$433 ( \4109 , \4010 , \4061 );
mand \mul_7_15/U$388 ( \4110 , \2955_A[8] , \2990_B[12] );
mand \mul_7_15/U$341 ( \4111 , \4109 , \4110 );
mxor \mul_7_15/U$342 ( \4112 , \4109 , \4110 );
mxor \mul_7_15/U$438 ( \4113 , \4014 , \4059 );
mand \mul_7_15/U$389 ( \4114 , \2959_A[7] , \2990_B[12] );
mand \mul_7_15/U$346 ( \4115 , \4113 , \4114 );
mxor \mul_7_15/U$347 ( \4116 , \4113 , \4114 );
mxor \mul_7_15/U$443 ( \4117 , \4018 , \4057 );
mand \mul_7_15/U$390 ( \4118 , \2963_A[6] , \2990_B[12] );
mand \mul_7_15/U$351 ( \4119 , \4117 , \4118 );
mxor \mul_7_15/U$352 ( \4120 , \4117 , \4118 );
mxor \mul_7_15/U$448 ( \4121 , \4022 , \4055 );
mand \mul_7_15/U$391 ( \4122 , \2967_A[5] , \2990_B[12] );
mand \mul_7_15/U$356 ( \4123 , \4121 , \4122 );
mxor \mul_7_15/U$357 ( \4124 , \4121 , \4122 );
mxor \mul_7_15/U$453 ( \4125 , \4026 , \4053 );
mand \mul_7_15/U$392 ( \4126 , \2971_A[4] , \2990_B[12] );
mand \mul_7_15/U$361 ( \4127 , \4125 , \4126 );
mxor \mul_7_15/U$362 ( \4128 , \4125 , \4126 );
mxor \mul_7_15/U$458 ( \4129 , \4030 , \4051 );
mand \mul_7_15/U$393 ( \4130 , \2975_A[3] , \2990_B[12] );
mand \mul_7_15/U$366 ( \4131 , \4129 , \4130 );
mxor \mul_7_15/U$367 ( \4132 , \4129 , \4130 );
mxor \mul_7_15/U$463 ( \4133 , \4034 , \4049 );
mand \mul_7_15/U$394 ( \4134 , \2979_A[2] , \2990_B[12] );
mand \mul_7_15/U$371 ( \4135 , \4133 , \4134 );
mxor \mul_7_15/U$372 ( \4136 , \4133 , \4134 );
mxor \mul_7_15/U$468 ( \4137 , \4038 , \4047 );
mand \mul_7_15/U$395 ( \4138 , \2983_A[1] , \2990_B[12] );
mand \mul_7_15/U$376 ( \4139 , \4137 , \4138 );
mxor \mul_7_15/U$377 ( \4140 , \4137 , \4138 );
mxor \mul_7_15/U$473 ( \4141 , \4042 , \4045 );
mand \mul_7_15/U$396 ( \4142 , \2986_A[0] , \2990_B[12] );
mand \mul_7_15/U$378 ( \4143 , \4141 , \4142 );
mand \mul_7_15/U$375 ( \4144 , \4140 , \4143 );
mor \mul_7_15/U$373 ( \4145 , \4139 , \4144 );
mand \mul_7_15/U$370 ( \4146 , \4136 , \4145 );
mor \mul_7_15/U$368 ( \4147 , \4135 , \4146 );
mand \mul_7_15/U$365 ( \4148 , \4132 , \4147 );
mor \mul_7_15/U$363 ( \4149 , \4131 , \4148 );
mand \mul_7_15/U$360 ( \4150 , \4128 , \4149 );
mor \mul_7_15/U$358 ( \4151 , \4127 , \4150 );
mand \mul_7_15/U$355 ( \4152 , \4124 , \4151 );
mor \mul_7_15/U$353 ( \4153 , \4123 , \4152 );
mand \mul_7_15/U$350 ( \4154 , \4120 , \4153 );
mor \mul_7_15/U$348 ( \4155 , \4119 , \4154 );
mand \mul_7_15/U$345 ( \4156 , \4116 , \4155 );
mor \mul_7_15/U$343 ( \4157 , \4115 , \4156 );
mand \mul_7_15/U$340 ( \4158 , \4112 , \4157 );
mor \mul_7_15/U$338 ( \4159 , \4111 , \4158 );
mand \mul_7_15/U$335 ( \4160 , \4108 , \4159 );
mor \mul_7_15/U$333 ( \4161 , \4107 , \4160 );
mand \mul_7_15/U$330 ( \4162 , \4104 , \4161 );
mor \mul_7_15/U$328 ( \4163 , \4103 , \4162 );
mand \mul_7_15/U$325 ( \4164 , \4100 , \4163 );
mor \mul_7_15/U$323 ( \4165 , \4099 , \4164 );
mand \mul_7_15/U$320 ( \4166 , \4096 , \4165 );
mor \mul_7_15/U$318 ( \4167 , \4095 , \4166 );
mand \mul_7_15/U$315 ( \4168 , \4092 , \4167 );
mor \mul_7_15/U$313 ( \4169 , \4091 , \4168 );
mand \mul_7_15/U$310 ( \4170 , \4088 , \4169 );
mor \mul_7_15/U$308 ( \4171 , \4087 , \4170 );
mand \mul_7_15/U$305 ( \4172 , \4084 , \4171 );
mor \mul_7_15/U$303 ( \4173 , \4083 , \4172 );
mand \mul_7_15/U$300 ( \4174 , \4080 , \4173 );
mor \mul_7_15/U$298 ( \4175 , \4079 , \4174 );
mand \mul_7_15/U$281 ( \4176 , \2923_A[16] , \2989_B[13] );
mand \mul_7_15/U$202 ( \4177 , \4175 , \4176 );
mxor \mul_7_15/U$203 ( \4178 , \4175 , \4176 );
mxor \mul_7_15/U$299 ( \4179 , \4080 , \4173 );
mand \mul_7_15/U$282 ( \4180 , \2927_A[15] , \2989_B[13] );
mand \mul_7_15/U$207 ( \4181 , \4179 , \4180 );
mxor \mul_7_15/U$208 ( \4182 , \4179 , \4180 );
mxor \mul_7_15/U$304 ( \4183 , \4084 , \4171 );
mand \mul_7_15/U$283 ( \4184 , \2931_A[14] , \2989_B[13] );
mand \mul_7_15/U$212 ( \4185 , \4183 , \4184 );
mxor \mul_7_15/U$213 ( \4186 , \4183 , \4184 );
mxor \mul_7_15/U$309 ( \4187 , \4088 , \4169 );
mand \mul_7_15/U$284 ( \4188 , \2935_A[13] , \2989_B[13] );
mand \mul_7_15/U$217 ( \4189 , \4187 , \4188 );
mxor \mul_7_15/U$218 ( \4190 , \4187 , \4188 );
mxor \mul_7_15/U$314 ( \4191 , \4092 , \4167 );
mand \mul_7_15/U$285 ( \4192 , \2939_A[12] , \2989_B[13] );
mand \mul_7_15/U$222 ( \4193 , \4191 , \4192 );
mxor \mul_7_15/U$223 ( \4194 , \4191 , \4192 );
mxor \mul_7_15/U$319 ( \4195 , \4096 , \4165 );
mand \mul_7_15/U$286 ( \4196 , \2943_A[11] , \2989_B[13] );
mand \mul_7_15/U$227 ( \4197 , \4195 , \4196 );
mxor \mul_7_15/U$228 ( \4198 , \4195 , \4196 );
mxor \mul_7_15/U$324 ( \4199 , \4100 , \4163 );
mand \mul_7_15/U$287 ( \4200 , \2947_A[10] , \2989_B[13] );
mand \mul_7_15/U$232 ( \4201 , \4199 , \4200 );
mxor \mul_7_15/U$233 ( \4202 , \4199 , \4200 );
mxor \mul_7_15/U$329 ( \4203 , \4104 , \4161 );
mand \mul_7_15/U$288 ( \4204 , \2951_A[9] , \2989_B[13] );
mand \mul_7_15/U$237 ( \4205 , \4203 , \4204 );
mxor \mul_7_15/U$238 ( \4206 , \4203 , \4204 );
mxor \mul_7_15/U$334 ( \4207 , \4108 , \4159 );
mand \mul_7_15/U$289 ( \4208 , \2955_A[8] , \2989_B[13] );
mand \mul_7_15/U$242 ( \4209 , \4207 , \4208 );
mxor \mul_7_15/U$243 ( \4210 , \4207 , \4208 );
mxor \mul_7_15/U$339 ( \4211 , \4112 , \4157 );
mand \mul_7_15/U$290 ( \4212 , \2959_A[7] , \2989_B[13] );
mand \mul_7_15/U$247 ( \4213 , \4211 , \4212 );
mxor \mul_7_15/U$248 ( \4214 , \4211 , \4212 );
mxor \mul_7_15/U$344 ( \4215 , \4116 , \4155 );
mand \mul_7_15/U$291 ( \4216 , \2963_A[6] , \2989_B[13] );
mand \mul_7_15/U$252 ( \4217 , \4215 , \4216 );
mxor \mul_7_15/U$253 ( \4218 , \4215 , \4216 );
mxor \mul_7_15/U$349 ( \4219 , \4120 , \4153 );
mand \mul_7_15/U$292 ( \4220 , \2967_A[5] , \2989_B[13] );
mand \mul_7_15/U$257 ( \4221 , \4219 , \4220 );
mxor \mul_7_15/U$258 ( \4222 , \4219 , \4220 );
mxor \mul_7_15/U$354 ( \4223 , \4124 , \4151 );
mand \mul_7_15/U$293 ( \4224 , \2971_A[4] , \2989_B[13] );
mand \mul_7_15/U$262 ( \4225 , \4223 , \4224 );
mxor \mul_7_15/U$263 ( \4226 , \4223 , \4224 );
mxor \mul_7_15/U$359 ( \4227 , \4128 , \4149 );
mand \mul_7_15/U$294 ( \4228 , \2975_A[3] , \2989_B[13] );
mand \mul_7_15/U$267 ( \4229 , \4227 , \4228 );
mxor \mul_7_15/U$268 ( \4230 , \4227 , \4228 );
mxor \mul_7_15/U$364 ( \4231 , \4132 , \4147 );
mand \mul_7_15/U$295 ( \4232 , \2979_A[2] , \2989_B[13] );
mand \mul_7_15/U$272 ( \4233 , \4231 , \4232 );
mxor \mul_7_15/U$273 ( \4234 , \4231 , \4232 );
mxor \mul_7_15/U$369 ( \4235 , \4136 , \4145 );
mand \mul_7_15/U$296 ( \4236 , \2983_A[1] , \2989_B[13] );
mand \mul_7_15/U$277 ( \4237 , \4235 , \4236 );
mxor \mul_7_15/U$278 ( \4238 , \4235 , \4236 );
mxor \mul_7_15/U$374 ( \4239 , \4140 , \4143 );
mand \mul_7_15/U$297 ( \4240 , \2986_A[0] , \2989_B[13] );
mand \mul_7_15/U$279 ( \4241 , \4239 , \4240 );
mand \mul_7_15/U$276 ( \4242 , \4238 , \4241 );
mor \mul_7_15/U$274 ( \4243 , \4237 , \4242 );
mand \mul_7_15/U$271 ( \4244 , \4234 , \4243 );
mor \mul_7_15/U$269 ( \4245 , \4233 , \4244 );
mand \mul_7_15/U$266 ( \4246 , \4230 , \4245 );
mor \mul_7_15/U$264 ( \4247 , \4229 , \4246 );
mand \mul_7_15/U$261 ( \4248 , \4226 , \4247 );
mor \mul_7_15/U$259 ( \4249 , \4225 , \4248 );
mand \mul_7_15/U$256 ( \4250 , \4222 , \4249 );
mor \mul_7_15/U$254 ( \4251 , \4221 , \4250 );
mand \mul_7_15/U$251 ( \4252 , \4218 , \4251 );
mor \mul_7_15/U$249 ( \4253 , \4217 , \4252 );
mand \mul_7_15/U$246 ( \4254 , \4214 , \4253 );
mor \mul_7_15/U$244 ( \4255 , \4213 , \4254 );
mand \mul_7_15/U$241 ( \4256 , \4210 , \4255 );
mor \mul_7_15/U$239 ( \4257 , \4209 , \4256 );
mand \mul_7_15/U$236 ( \4258 , \4206 , \4257 );
mor \mul_7_15/U$234 ( \4259 , \4205 , \4258 );
mand \mul_7_15/U$231 ( \4260 , \4202 , \4259 );
mor \mul_7_15/U$229 ( \4261 , \4201 , \4260 );
mand \mul_7_15/U$226 ( \4262 , \4198 , \4261 );
mor \mul_7_15/U$224 ( \4263 , \4197 , \4262 );
mand \mul_7_15/U$221 ( \4264 , \4194 , \4263 );
mor \mul_7_15/U$219 ( \4265 , \4193 , \4264 );
mand \mul_7_15/U$216 ( \4266 , \4190 , \4265 );
mor \mul_7_15/U$214 ( \4267 , \4189 , \4266 );
mand \mul_7_15/U$211 ( \4268 , \4186 , \4267 );
mor \mul_7_15/U$209 ( \4269 , \4185 , \4268 );
mand \mul_7_15/U$206 ( \4270 , \4182 , \4269 );
mor \mul_7_15/U$204 ( \4271 , \4181 , \4270 );
mand \mul_7_15/U$201 ( \4272 , \4178 , \4271 );
mor \mul_7_15/U$199 ( \4273 , \4177 , \4272 );
mand \mul_7_15/U$182 ( \4274 , \2923_A[16] , \2988_B[14] );
mand \mul_7_15/U$103 ( \4275 , \4273 , \4274 );
mxor \mul_7_15/U$104 ( \4276 , \4273 , \4274 );
mxor \mul_7_15/U$200 ( \4277 , \4178 , \4271 );
mand \mul_7_15/U$183 ( \4278 , \2927_A[15] , \2988_B[14] );
mand \mul_7_15/U$108 ( \4279 , \4277 , \4278 );
mxor \mul_7_15/U$109 ( \4280 , \4277 , \4278 );
mxor \mul_7_15/U$205 ( \4281 , \4182 , \4269 );
mand \mul_7_15/U$184 ( \4282 , \2931_A[14] , \2988_B[14] );
mand \mul_7_15/U$113 ( \4283 , \4281 , \4282 );
mxor \mul_7_15/U$114 ( \4284 , \4281 , \4282 );
mxor \mul_7_15/U$210 ( \4285 , \4186 , \4267 );
mand \mul_7_15/U$185 ( \4286 , \2935_A[13] , \2988_B[14] );
mand \mul_7_15/U$118 ( \4287 , \4285 , \4286 );
mxor \mul_7_15/U$119 ( \4288 , \4285 , \4286 );
mxor \mul_7_15/U$215 ( \4289 , \4190 , \4265 );
mand \mul_7_15/U$186 ( \4290 , \2939_A[12] , \2988_B[14] );
mand \mul_7_15/U$123 ( \4291 , \4289 , \4290 );
mxor \mul_7_15/U$124 ( \4292 , \4289 , \4290 );
mxor \mul_7_15/U$220 ( \4293 , \4194 , \4263 );
mand \mul_7_15/U$187 ( \4294 , \2943_A[11] , \2988_B[14] );
mand \mul_7_15/U$128 ( \4295 , \4293 , \4294 );
mxor \mul_7_15/U$129 ( \4296 , \4293 , \4294 );
mxor \mul_7_15/U$225 ( \4297 , \4198 , \4261 );
mand \mul_7_15/U$188 ( \4298 , \2947_A[10] , \2988_B[14] );
mand \mul_7_15/U$133 ( \4299 , \4297 , \4298 );
mxor \mul_7_15/U$134 ( \4300 , \4297 , \4298 );
mxor \mul_7_15/U$230 ( \4301 , \4202 , \4259 );
mand \mul_7_15/U$189 ( \4302 , \2951_A[9] , \2988_B[14] );
mand \mul_7_15/U$138 ( \4303 , \4301 , \4302 );
mxor \mul_7_15/U$139 ( \4304 , \4301 , \4302 );
mxor \mul_7_15/U$235 ( \4305 , \4206 , \4257 );
mand \mul_7_15/U$190 ( \4306 , \2955_A[8] , \2988_B[14] );
mand \mul_7_15/U$143 ( \4307 , \4305 , \4306 );
mxor \mul_7_15/U$144 ( \4308 , \4305 , \4306 );
mxor \mul_7_15/U$240 ( \4309 , \4210 , \4255 );
mand \mul_7_15/U$191 ( \4310 , \2959_A[7] , \2988_B[14] );
mand \mul_7_15/U$148 ( \4311 , \4309 , \4310 );
mxor \mul_7_15/U$149 ( \4312 , \4309 , \4310 );
mxor \mul_7_15/U$245 ( \4313 , \4214 , \4253 );
mand \mul_7_15/U$192 ( \4314 , \2963_A[6] , \2988_B[14] );
mand \mul_7_15/U$153 ( \4315 , \4313 , \4314 );
mxor \mul_7_15/U$154 ( \4316 , \4313 , \4314 );
mxor \mul_7_15/U$250 ( \4317 , \4218 , \4251 );
mand \mul_7_15/U$193 ( \4318 , \2967_A[5] , \2988_B[14] );
mand \mul_7_15/U$158 ( \4319 , \4317 , \4318 );
mxor \mul_7_15/U$159 ( \4320 , \4317 , \4318 );
mxor \mul_7_15/U$255 ( \4321 , \4222 , \4249 );
mand \mul_7_15/U$194 ( \4322 , \2971_A[4] , \2988_B[14] );
mand \mul_7_15/U$163 ( \4323 , \4321 , \4322 );
mxor \mul_7_15/U$164 ( \4324 , \4321 , \4322 );
mxor \mul_7_15/U$260 ( \4325 , \4226 , \4247 );
mand \mul_7_15/U$195 ( \4326 , \2975_A[3] , \2988_B[14] );
mand \mul_7_15/U$168 ( \4327 , \4325 , \4326 );
mxor \mul_7_15/U$169 ( \4328 , \4325 , \4326 );
mxor \mul_7_15/U$265 ( \4329 , \4230 , \4245 );
mand \mul_7_15/U$196 ( \4330 , \2979_A[2] , \2988_B[14] );
mand \mul_7_15/U$173 ( \4331 , \4329 , \4330 );
mxor \mul_7_15/U$174 ( \4332 , \4329 , \4330 );
mxor \mul_7_15/U$270 ( \4333 , \4234 , \4243 );
mand \mul_7_15/U$197 ( \4334 , \2983_A[1] , \2988_B[14] );
mand \mul_7_15/U$178 ( \4335 , \4333 , \4334 );
mxor \mul_7_15/U$179 ( \4336 , \4333 , \4334 );
mxor \mul_7_15/U$275 ( \4337 , \4238 , \4241 );
mand \mul_7_15/U$198 ( \4338 , \2986_A[0] , \2988_B[14] );
mand \mul_7_15/U$180 ( \4339 , \4337 , \4338 );
mand \mul_7_15/U$177 ( \4340 , \4336 , \4339 );
mor \mul_7_15/U$175 ( \4341 , \4335 , \4340 );
mand \mul_7_15/U$172 ( \4342 , \4332 , \4341 );
mor \mul_7_15/U$170 ( \4343 , \4331 , \4342 );
mand \mul_7_15/U$167 ( \4344 , \4328 , \4343 );
mor \mul_7_15/U$165 ( \4345 , \4327 , \4344 );
mand \mul_7_15/U$162 ( \4346 , \4324 , \4345 );
mor \mul_7_15/U$160 ( \4347 , \4323 , \4346 );
mand \mul_7_15/U$157 ( \4348 , \4320 , \4347 );
mor \mul_7_15/U$155 ( \4349 , \4319 , \4348 );
mand \mul_7_15/U$152 ( \4350 , \4316 , \4349 );
mor \mul_7_15/U$150 ( \4351 , \4315 , \4350 );
mand \mul_7_15/U$147 ( \4352 , \4312 , \4351 );
mor \mul_7_15/U$145 ( \4353 , \4311 , \4352 );
mand \mul_7_15/U$142 ( \4354 , \4308 , \4353 );
mor \mul_7_15/U$140 ( \4355 , \4307 , \4354 );
mand \mul_7_15/U$137 ( \4356 , \4304 , \4355 );
mor \mul_7_15/U$135 ( \4357 , \4303 , \4356 );
mand \mul_7_15/U$132 ( \4358 , \4300 , \4357 );
mor \mul_7_15/U$130 ( \4359 , \4299 , \4358 );
mand \mul_7_15/U$127 ( \4360 , \4296 , \4359 );
mor \mul_7_15/U$125 ( \4361 , \4295 , \4360 );
mand \mul_7_15/U$122 ( \4362 , \4292 , \4361 );
mor \mul_7_15/U$120 ( \4363 , \4291 , \4362 );
mand \mul_7_15/U$117 ( \4364 , \4288 , \4363 );
mor \mul_7_15/U$115 ( \4365 , \4287 , \4364 );
mand \mul_7_15/U$112 ( \4366 , \4284 , \4365 );
mor \mul_7_15/U$110 ( \4367 , \4283 , \4366 );
mand \mul_7_15/U$107 ( \4368 , \4280 , \4367 );
mor \mul_7_15/U$105 ( \4369 , \4279 , \4368 );
mand \mul_7_15/U$102 ( \4370 , \4276 , \4369 );
mor \mul_7_15/U$100 ( \4371 , \4275 , \4370 );
mand \mul_7_15/U$83 ( \4372 , \2923_A[16] , \2987_B[15] );
mxor \mul_7_15/U$5 ( \4373 , \4371 , \4372 );
mxor \mul_7_15/U$101 ( \4374 , \4276 , \4369 );
mand \mul_7_15/U$84 ( \4375 , \2927_A[15] , \2987_B[15] );
mand \mul_7_15/U$9 ( \4376 , \4374 , \4375 );
mxor \mul_7_15/U$10 ( \4377 , \4374 , \4375 );
mxor \mul_7_15/U$106 ( \4378 , \4280 , \4367 );
mand \mul_7_15/U$85 ( \4379 , \2931_A[14] , \2987_B[15] );
mand \mul_7_15/U$14 ( \4380 , \4378 , \4379 );
mxor \mul_7_15/U$15 ( \4381 , \4378 , \4379 );
mxor \mul_7_15/U$111 ( \4382 , \4284 , \4365 );
mand \mul_7_15/U$86 ( \4383 , \2935_A[13] , \2987_B[15] );
mand \mul_7_15/U$19 ( \4384 , \4382 , \4383 );
mxor \mul_7_15/U$20 ( \4385 , \4382 , \4383 );
mxor \mul_7_15/U$116 ( \4386 , \4288 , \4363 );
mand \mul_7_15/U$87 ( \4387 , \2939_A[12] , \2987_B[15] );
mand \mul_7_15/U$24 ( \4388 , \4386 , \4387 );
mxor \mul_7_15/U$25 ( \4389 , \4386 , \4387 );
mxor \mul_7_15/U$121 ( \4390 , \4292 , \4361 );
mand \mul_7_15/U$88 ( \4391 , \2943_A[11] , \2987_B[15] );
mand \mul_7_15/U$29 ( \4392 , \4390 , \4391 );
mxor \mul_7_15/U$30 ( \4393 , \4390 , \4391 );
mxor \mul_7_15/U$126 ( \4394 , \4296 , \4359 );
mand \mul_7_15/U$89 ( \4395 , \2947_A[10] , \2987_B[15] );
mand \mul_7_15/U$34 ( \4396 , \4394 , \4395 );
mxor \mul_7_15/U$35 ( \4397 , \4394 , \4395 );
mxor \mul_7_15/U$131 ( \4398 , \4300 , \4357 );
mand \mul_7_15/U$90 ( \4399 , \2951_A[9] , \2987_B[15] );
mand \mul_7_15/U$39 ( \4400 , \4398 , \4399 );
mxor \mul_7_15/U$40 ( \4401 , \4398 , \4399 );
mxor \mul_7_15/U$136 ( \4402 , \4304 , \4355 );
mand \mul_7_15/U$91 ( \4403 , \2955_A[8] , \2987_B[15] );
mand \mul_7_15/U$44 ( \4404 , \4402 , \4403 );
mxor \mul_7_15/U$45 ( \4405 , \4402 , \4403 );
mxor \mul_7_15/U$141 ( \4406 , \4308 , \4353 );
mand \mul_7_15/U$92 ( \4407 , \2959_A[7] , \2987_B[15] );
mand \mul_7_15/U$49 ( \4408 , \4406 , \4407 );
mxor \mul_7_15/U$50 ( \4409 , \4406 , \4407 );
mxor \mul_7_15/U$146 ( \4410 , \4312 , \4351 );
mand \mul_7_15/U$93 ( \4411 , \2963_A[6] , \2987_B[15] );
mand \mul_7_15/U$54 ( \4412 , \4410 , \4411 );
mxor \mul_7_15/U$55 ( \4413 , \4410 , \4411 );
mxor \mul_7_15/U$151 ( \4414 , \4316 , \4349 );
mand \mul_7_15/U$94 ( \4415 , \2967_A[5] , \2987_B[15] );
mand \mul_7_15/U$59 ( \4416 , \4414 , \4415 );
mxor \mul_7_15/U$60 ( \4417 , \4414 , \4415 );
mxor \mul_7_15/U$156 ( \4418 , \4320 , \4347 );
mand \mul_7_15/U$95 ( \4419 , \2971_A[4] , \2987_B[15] );
mand \mul_7_15/U$64 ( \4420 , \4418 , \4419 );
mxor \mul_7_15/U$65 ( \4421 , \4418 , \4419 );
mxor \mul_7_15/U$161 ( \4422 , \4324 , \4345 );
mand \mul_7_15/U$96 ( \4423 , \2975_A[3] , \2987_B[15] );
mand \mul_7_15/U$69 ( \4424 , \4422 , \4423 );
mxor \mul_7_15/U$70 ( \4425 , \4422 , \4423 );
mxor \mul_7_15/U$166 ( \4426 , \4328 , \4343 );
mand \mul_7_15/U$97 ( \4427 , \2979_A[2] , \2987_B[15] );
mand \mul_7_15/U$74 ( \4428 , \4426 , \4427 );
mxor \mul_7_15/U$75 ( \4429 , \4426 , \4427 );
mxor \mul_7_15/U$171 ( \4430 , \4332 , \4341 );
mand \mul_7_15/U$98 ( \4431 , \2983_A[1] , \2987_B[15] );
mand \mul_7_15/U$79 ( \4432 , \4430 , \4431 );
mxor \mul_7_15/U$80 ( \4433 , \4430 , \4431 );
mxor \mul_7_15/U$176 ( \4434 , \4336 , \4339 );
mand \mul_7_15/U$99 ( \4435 , \2986_A[0] , \2987_B[15] );
mand \mul_7_15/U$81 ( \4436 , \4434 , \4435 );
mand \mul_7_15/U$78 ( \4437 , \4433 , \4436 );
mor \mul_7_15/U$76 ( \4438 , \4432 , \4437 );
mand \mul_7_15/U$73 ( \4439 , \4429 , \4438 );
mor \mul_7_15/U$71 ( \4440 , \4428 , \4439 );
mand \mul_7_15/U$68 ( \4441 , \4425 , \4440 );
mor \mul_7_15/U$66 ( \4442 , \4424 , \4441 );
mand \mul_7_15/U$63 ( \4443 , \4421 , \4442 );
mor \mul_7_15/U$61 ( \4444 , \4420 , \4443 );
mand \mul_7_15/U$58 ( \4445 , \4417 , \4444 );
mor \mul_7_15/U$56 ( \4446 , \4416 , \4445 );
mand \mul_7_15/U$53 ( \4447 , \4413 , \4446 );
mor \mul_7_15/U$51 ( \4448 , \4412 , \4447 );
mand \mul_7_15/U$48 ( \4449 , \4409 , \4448 );
mor \mul_7_15/U$46 ( \4450 , \4408 , \4449 );
mand \mul_7_15/U$43 ( \4451 , \4405 , \4450 );
mor \mul_7_15/U$41 ( \4452 , \4404 , \4451 );
mand \mul_7_15/U$38 ( \4453 , \4401 , \4452 );
mor \mul_7_15/U$36 ( \4454 , \4400 , \4453 );
mand \mul_7_15/U$33 ( \4455 , \4397 , \4454 );
mor \mul_7_15/U$31 ( \4456 , \4396 , \4455 );
mand \mul_7_15/U$28 ( \4457 , \4393 , \4456 );
mor \mul_7_15/U$26 ( \4458 , \4392 , \4457 );
mand \mul_7_15/U$23 ( \4459 , \4389 , \4458 );
mor \mul_7_15/U$21 ( \4460 , \4388 , \4459 );
mand \mul_7_15/U$18 ( \4461 , \4385 , \4460 );
mor \mul_7_15/U$16 ( \4462 , \4384 , \4461 );
mand \mul_7_15/U$13 ( \4463 , \4381 , \4462 );
mor \mul_7_15/U$11 ( \4464 , \4380 , \4463 );
mand \mul_7_15/U$8 ( \4465 , \4377 , \4464 );
mor \mul_7_15/U$6 ( \4466 , \4376 , \4465 );
mxor \mul_7_15/U$2 ( \4467 , \4373 , \4466 );
mbuf \mul_7_15/Z[31] ( \4468_Z[31] , \4467 );
mxor \mul_7_15/U$7 ( \4469 , \4377 , \4464 );
mbuf \mul_7_15/Z[30] ( \4470_Z[30] , \4469 );
mxor \mul_7_15/U$12 ( \4471 , \4381 , \4462 );
mbuf \mul_7_15/Z[29] ( \4472_Z[29] , \4471 );
mxor \mul_7_15/U$17 ( \4473 , \4385 , \4460 );
mbuf \mul_7_15/Z[28] ( \4474_Z[28] , \4473 );
mxor \mul_7_15/U$22 ( \4475 , \4389 , \4458 );
mbuf \mul_7_15/Z[27] ( \4476_Z[27] , \4475 );
mxor \mul_7_15/U$27 ( \4477 , \4393 , \4456 );
mbuf \mul_7_15/Z[26] ( \4478_Z[26] , \4477 );
mxor \mul_7_15/U$32 ( \4479 , \4397 , \4454 );
mbuf \mul_7_15/Z[25] ( \4480_Z[25] , \4479 );
mxor \mul_7_15/U$37 ( \4481 , \4401 , \4452 );
mbuf \mul_7_15/Z[24] ( \4482_Z[24] , \4481 );
mxor \mul_7_15/U$42 ( \4483 , \4405 , \4450 );
mbuf \mul_7_15/Z[23] ( \4484_Z[23] , \4483 );
mxor \mul_7_15/U$47 ( \4485 , \4409 , \4448 );
mbuf \mul_7_15/Z[22] ( \4486_Z[22] , \4485 );
mxor \mul_7_15/U$52 ( \4487 , \4413 , \4446 );
mbuf \mul_7_15/Z[21] ( \4488_Z[21] , \4487 );
mxor \mul_7_15/U$57 ( \4489 , \4417 , \4444 );
mbuf \mul_7_15/Z[20] ( \4490_Z[20] , \4489 );
mxor \mul_7_15/U$62 ( \4491 , \4421 , \4442 );
mbuf \mul_7_15/Z[19] ( \4492_Z[19] , \4491 );
mxor \mul_7_15/U$67 ( \4493 , \4425 , \4440 );
mbuf \mul_7_15/Z[18] ( \4494_Z[18] , \4493 );
mxor \mul_7_15/U$72 ( \4495 , \4429 , \4438 );
mbuf \mul_7_15/Z[17] ( \4496_Z[17] , \4495 );
mxor \mul_7_15/U$77 ( \4497 , \4433 , \4436 );
mbuf \mul_7_15/Z[16] ( \4498_Z[16] , \4497 );
mxor \mul_7_15/U$82 ( \4499 , \4434 , \4435 );
mbuf \mul_7_15/Z[15] ( \4500_Z[15] , \4499 );
mxor \mul_7_15/U$181 ( \4501 , \4337 , \4338 );
mbuf \mul_7_15/Z[14] ( \4502_Z[14] , \4501 );
mxor \mul_7_15/U$280 ( \4503 , \4239 , \4240 );
mbuf \mul_7_15/Z[13] ( \4504_Z[13] , \4503 );
mxor \mul_7_15/U$379 ( \4505 , \4141 , \4142 );
mbuf \mul_7_15/Z[12] ( \4506_Z[12] , \4505 );
mxor \mul_7_15/U$478 ( \4507 , \4043 , \4044 );
mbuf \mul_7_15/Z[11] ( \4508_Z[11] , \4507 );
mxor \mul_7_15/U$577 ( \4509 , \3945 , \3946 );
mbuf \mul_7_15/Z[10] ( \4510_Z[10] , \4509 );
mxor \mul_7_15/U$676 ( \4511 , \3847 , \3848 );
mbuf \mul_7_15/Z[9] ( \4512_Z[9] , \4511 );
mxor \mul_7_15/U$775 ( \4513 , \3749 , \3750 );
mbuf \mul_7_15/Z[8] ( \4514_Z[8] , \4513 );
mxor \mul_7_15/U$874 ( \4515 , \3651 , \3652 );
mbuf \mul_7_15/Z[7] ( \4516_Z[7] , \4515 );
mxor \mul_7_15/U$973 ( \4517 , \3553 , \3554 );
mbuf \mul_7_15/Z[6] ( \4518_Z[6] , \4517 );
mxor \mul_7_15/U$1072 ( \4519 , \3455 , \3456 );
mbuf \mul_7_15/Z[5] ( \4520_Z[5] , \4519 );
mxor \mul_7_15/U$1171 ( \4521 , \3357 , \3358 );
mbuf \mul_7_15/Z[4] ( \4522_Z[4] , \4521 );
mxor \mul_7_15/U$1270 ( \4523 , \3259 , \3260 );
mbuf \mul_7_15/Z[3] ( \4524_Z[3] , \4523 );
mxor \mul_7_15/U$1369 ( \4525 , \3161 , \3162 );
mbuf \mul_7_15/Z[2] ( \4526_Z[2] , \4525 );
mxor \mul_7_15/U$1465 ( \4527 , \3064 , \3065 );
mbuf \mul_7_15/Z[1] ( \4528_Z[1] , \4527 );
mand \mul_7_15/U$1499 ( \4529 , \2986_A[0] , \3002_B[0] );
mbuf \mul_7_15/Z[0] ( \4530_Z[0] , \4529 );
endmodule


//
// Conformal-LEC Version 19.20-d255 (16-Apr-2020)
//
module top(\a[15] ,\a[14] ,\a[13] ,\a[12] ,\a[11] ,\a[10] ,\a[9] ,\a[8] ,\a[7] ,
        \a[6] ,\a[5] ,\a[4] ,\a[3] ,\a[2] ,\a[1] ,\a[0] ,\b[15] ,\b[14] ,\b[13] ,
        \b[12] ,\b[11] ,\b[10] ,\b[9] ,\b[8] ,\b[7] ,\b[6] ,\b[5] ,\b[4] ,\b[3] ,
        \b[2] ,\b[1] ,\b[0] ,\c[15] ,\c[14] ,\c[13] ,\c[12] ,\c[11] ,\c[10] ,\c[9] ,
        \c[8] ,\c[7] ,\c[6] ,\c[5] ,\c[4] ,\c[3] ,\c[2] ,\c[1] ,\c[0] ,\d[15] ,
        \d[14] ,\d[13] ,\d[12] ,\d[11] ,\d[10] ,\d[9] ,\d[8] ,\d[7] ,\d[6] ,\d[5] ,
        \d[4] ,\d[3] ,\d[2] ,\d[1] ,\d[0] ,\o[31] ,\o[30] ,\o[29] ,\o[28] ,\o[27] ,
        \o[26] ,\o[25] ,\o[24] ,\o[23] ,\o[22] ,\o[21] ,\o[20] ,\o[19] ,\o[18] ,\o[17] ,
        \o[16] ,\o[15] ,\o[14] ,\o[13] ,\o[12] ,\o[11] ,\o[10] ,\o[9] ,\o[8] ,\o[7] ,
        \o[6] ,\o[5] ,\o[4] ,\o[3] ,\o[2] ,\o[1] ,\o[0] );
input [1:0] \a[15] ,\a[14] ,\a[13] ,\a[12] ,\a[11] ,\a[10] ,\a[9] ,\a[8] ,\a[7] ,        \a[6] ,\a[5] ,\a[4] ,\a[3] ,\a[2] ,\a[1] ,\a[0] ,\b[15] ,\b[14] ,\b[13] ,        \b[12] ,\b[11] ,\b[10] ,\b[9] ,\b[8] ,\b[7] ,\b[6] ,\b[5] ,\b[4] ,\b[3] ,        \b[2] ,\b[1] ,\b[0] ,\c[15] ,\c[14] ,\c[13] ,\c[12] ,\c[11] ,\c[10] ,\c[9] ,        \c[8] ,\c[7] ,\c[6] ,\c[5] ,\c[4] ,\c[3] ,\c[2] ,\c[1] ,\c[0] ,\d[15] ,        \d[14] ,\d[13] ,\d[12] ,\d[11] ,\d[10] ,\d[9] ,\d[8] ,\d[7] ,\d[6] ,\d[5] ,        \d[4] ,\d[3] ,\d[2] ,\d[1] ,\d[0] ;
output [1:0] \o[31] ,\o[30] ,\o[29] ,\o[28] ,\o[27] ,\o[26] ,\o[25] ,\o[24] ,\o[23] ,        \o[22] ,\o[21] ,\o[20] ,\o[19] ,\o[18] ,\o[17] ,\o[16] ,\o[15] ,\o[14] ,\o[13] ,        \o[12] ,\o[11] ,\o[10] ,\o[9] ,\o[8] ,\o[7] ,\o[6] ,\o[5] ,\o[4] ,\o[3] ,        \o[2] ,\o[1] ,\o[0] ;

wire [1:0] \97_ZERO , \98_ONE , \99 , \100 , \101 , \102 , \103 , \104 , \105 ,         \106 , \107 , \108 , \109 , \110 , \111 , \112 , \113 , \114 , \115 ,         \116 , \117 , \118 , \119 , \120 , \121 , \122 , \123 , \124 , \125 ,         \126 , \127 , \128 , \129 , \130 , \131 , \132 , \133 , \134 , \135 ,         \136 , \137 , \138 , \139 , \140 , \141 , \142 , \143 , \144 , \145 ,         \146 , \147 , \148 , \149 , \150 , \151 , \152 , \153 , \154 , \155 ,         \156 , \157 , \158 , \159 , \160 , \161 , \162 , \163 , \164 , \165 ,         \166 , \167 , \168 , \169 , \170 , \171 , \172 , \173 , \174 , \175 ,         \176 , \177 , \178 , \179 , \180 , \181 , \182 , \183 , \184 , \185 ,         \186 , \187 , \188 , \189 , \190 , \191 , \192 , \193 , \194 , \195 ,         \196 , \197 , \198 , \199 , \200 , \201 , \202 , \203 , \204 , \205 ,         \206 , \207 , \208 , \209 , \210 , \211 , \212 , \213 , \214 , \215 ,         \216 , \217 , \218 , \219 , \220 , \221 , \222 , \223 , \224 , \225 ,         \226 , \227 , \228 , \229 , \230 , \231 , \232 , \233 , \234 , \235 ,         \236 , \237 , \238 , \239 , \240 , \241 , \242 , \243 , \244 , \245 ,         \246 , \247 , \248 , \249 , \250 , \251 , \252 , \253 , \254 , \255 ,         \256 , \257 , \258 , \259 , \260 , \261 , \262 , \263 , \264 , \265 ,         \266 , \267 , \268 , \269 , \270 , \271 , \272 , \273 , \274 , \275 ,         \276 , \277 , \278 , \279 , \280 , \281 , \282 , \283 , \284 , \285 ,         \286 , \287 , \288 , \289 , \290 , \291 , \292 , \293 , \294 , \295 ,         \296 , \297 , \298 , \299 , \300 , \301 , \302 , \303 , \304 , \305 ,         \306 , \307 , \308 , \309 , \310 , \311 , \312 , \313 , \314 , \315 ,         \316 , \317 , \318 , \319 , \320 , \321 , \322 , \323 , \324 , \325 ,         \326 , \327 , \328 , \329 , \330 , \331 , \332 , \333 , \334 , \335 ,         \336 , \337 , \338 , \339 , \340 , \341 , \342 , \343 , \344 , \345 ,         \346 , \347 , \348 , \349 , \350 , \351 , \352 , \353 , \354 , \355 ,         \356 , \357 , \358 , \359 , \360 , \361 , \362 , \363 , \364 , \365 ,         \366 , \367 , \368 , \369 , \370 , \371 , \372 , \373 , \374 , \375 ,         \376 , \377 , \378 , \379 , \380 , \381 , \382 , \383 , \384 , \385 ,         \386 , \387 , \388 , \389 , \390 , \391 , \392 , \393 , \394 , \395 ,         \396 , \397 , \398 , \399 , \400 , \401 , \402 , \403 , \404 , \405 ,         \406 , \407 , \408 , \409 , \410 , \411 , \412 , \413 , \414 , \415 ,         \416 , \417 , \418 , \419 , \420 , \421 , \422 , \423 , \424 , \425 ,         \426 , \427 , \428 , \429 , \430 , \431 , \432 , \433 , \434 , \435 ,         \436 , \437 , \438 , \439 , \440 , \441 , \442 , \443 , \444 , \445 ,         \446 , \447 , \448 , \449 , \450 , \451 , \452 , \453 , \454 , \455 ,         \456 , \457 , \458 , \459 , \460 , \461 , \462 , \463 , \464 , \465 ,         \466 , \467 , \468 , \469 , \470 , \471 , \472 , \473 , \474 , \475 ,         \476 , \477 , \478 , \479 , \480 , \481 , \482 , \483 , \484 , \485 ,         \486 , \487 , \488 , \489 , \490 , \491 , \492 , \493 , \494 , \495 ,         \496 , \497 , \498 , \499 , \500 , \501 , \502 , \503 , \504 , \505 ,         \506 , \507 , \508 , \509 , \510 , \511 , \512 , \513 , \514 , \515 ,         \516 , \517 , \518 , \519 , \520 , \521 , \522 , \523 , \524 , \525 ,         \526 , \527 , \528 , \529 , \530 , \531 , \532 , \533 , \534 , \535 ,         \536 , \537 , \538 , \539 , \540 , \541 , \542 , \543 , \544 , \545 ,         \546 , \547 , \548 , \549 , \550 , \551 , \552 , \553 , \554 , \555 ,         \556 , \557 , \558 , \559 , \560 , \561 , \562 , \563 , \564 , \565 ,         \566 , \567 , \568 , \569 , \570 , \571 , \572 , \573 , \574 , \575 ,         \576 , \577 , \578 , \579 , \580 , \581 , \582 , \583 , \584 , \585 ,         \586 , \587 , \588 , \589 , \590 , \591 , \592 , \593 , \594 , \595 ,         \596 , \597 , \598 , \599 , \600 , \601 , \602 , \603 , \604 , \605 ,         \606 , \607 , \608 , \609 , \610 , \611 , \612 , \613 , \614 , \615 ,         \616 , \617 , \618 , \619 , \620 , \621 , \622 , \623 , \624 , \625 ,         \626 , \627 , \628 , \629 , \630 , \631 , \632 , \633 , \634 , \635 ,         \636 , \637 , \638 , \639 , \640 , \641 , \642 , \643 , \644 , \645 ,         \646 , \647 , \648 , \649 , \650 , \651 , \652 , \653 , \654 , \655 ,         \656 , \657 , \658 , \659 , \660 , \661 , \662 , \663 , \664 , \665 ,         \666 , \667 , \668 , \669 , \670 , \671 , \672 , \673 , \674 , \675 ,         \676 , \677 , \678 , \679 , \680 , \681 , \682 , \683 , \684 , \685 ,         \686 , \687 , \688 , \689 , \690 , \691 , \692 , \693 , \694 , \695 ,         \696 , \697 , \698 , \699 , \700 , \701 , \702 , \703 , \704 , \705 ,         \706 , \707 , \708 , \709 , \710 , \711 , \712 , \713 , \714 , \715 ,         \716 , \717 , \718 , \719 , \720 , \721 , \722 , \723 , \724 , \725 ,         \726 , \727 , \728 , \729 , \730 , \731 , \732 , \733 , \734 , \735 ,         \736 , \737 , \738 , \739 , \740 , \741 , \742 , \743 , \744 , \745 ,         \746 , \747 , \748 , \749 , \750 , \751 , \752 , \753 , \754 , \755 ,         \756 , \757 , \758 , \759 , \760 , \761 , \762 , \763 , \764 , \765 ,         \766 , \767 , \768 , \769 , \770 , \771 , \772 , \773 , \774 , \775 ,         \776 , \777 , \778 , \779 , \780 , \781 , \782 , \783 , \784 , \785 ,         \786 , \787 , \788 , \789 , \790 , \791 , \792 , \793 , \794 , \795 ,         \796 , \797 , \798 , \799 , \800 , \801 , \802 , \803 , \804 , \805 ,         \806 , \807 , \808 , \809 , \810 , \811 , \812 , \813 , \814 , \815 ,         \816 , \817 , \818 , \819 , \820 , \821 , \822 , \823 , \824 , \825 ,         \826 , \827 , \828 , \829 , \830 , \831 , \832 , \833 , \834 , \835 ,         \836 , \837 , \838 , \839 , \840 , \841 , \842 , \843 , \844 , \845 ,         \846 , \847 , \848 , \849 , \850 , \851 , \852 , \853 , \854 , \855 ,         \856 , \857 , \858 , \859 , \860 , \861 , \862 , \863 , \864 , \865 ,         \866 , \867 , \868 , \869 , \870 , \871 , \872 , \873 , \874 , \875 ,         \876 , \877 , \878 , \879 , \880 , \881 , \882 , \883 , \884 , \885 ,         \886 , \887 , \888 , \889 , \890 , \891 , \892 , \893 , \894 , \895 ,         \896 , \897 , \898 , \899 , \900 , \901 , \902 , \903 , \904 , \905 ,         \906 , \907 , \908 , \909 , \910 , \911 , \912 , \913 , \914 , \915 ,         \916 , \917 , \918 , \919 , \920 , \921 , \922 , \923 , \924 , \925 ,         \926 , \927 , \928 , \929 , \930 , \931 , \932 , \933 , \934 , \935 ,         \936 , \937 , \938 , \939 , \940 , \941 , \942 , \943 , \944 , \945 ,         \946 , \947 , \948 , \949 , \950 , \951 , \952 , \953 , \954 , \955 ,         \956 , \957 , \958 , \959 , \960 , \961 , \962 , \963 , \964 , \965 ,         \966 , \967 , \968 , \969 , \970 , \971 , \972 , \973 , \974 , \975 ,         \976 , \977 , \978 , \979 , \980 , \981 , \982 , \983 , \984 , \985 ,         \986 , \987 , \988 , \989 , \990 , \991 , \992 , \993 , \994 , \995 ,         \996 , \997 , \998 , \999 , \1000 , \1001 , \1002 , \1003 , \1004 , \1005 ,         \1006 , \1007 , \1008 , \1009 , \1010 , \1011 , \1012 , \1013 , \1014 , \1015 ,         \1016 , \1017 , \1018 , \1019 , \1020 , \1021 , \1022 , \1023 , \1024 , \1025 ,         \1026 , \1027 , \1028 , \1029 , \1030 , \1031 , \1032 , \1033 , \1034 , \1035 ,         \1036 , \1037 , \1038 , \1039 , \1040 , \1041 , \1042 , \1043 , \1044 , \1045 ,         \1046 , \1047 , \1048 , \1049 , \1050 , \1051 , \1052 , \1053 , \1054 , \1055 ,         \1056 , \1057 , \1058 , \1059 , \1060 , \1061 , \1062 , \1063 , \1064 , \1065 ,         \1066 , \1067 , \1068 , \1069 , \1070 , \1071 , \1072 , \1073 , \1074 , \1075 ,         \1076 , \1077 , \1078 , \1079 , \1080 , \1081 , \1082 , \1083 , \1084 , \1085 ,         \1086 , \1087 , \1088 , \1089 , \1090 , \1091 , \1092 , \1093 , \1094 , \1095 ,         \1096 , \1097 , \1098 , \1099 , \1100 , \1101 , \1102 , \1103 , \1104 , \1105 ,         \1106 , \1107 , \1108 , \1109 , \1110 , \1111 , \1112 , \1113 , \1114 , \1115 ,         \1116 , \1117 , \1118 , \1119 , \1120 , \1121 , \1122 , \1123 , \1124 , \1125 ,         \1126 , \1127 , \1128 , \1129 , \1130 , \1131 , \1132 , \1133 , \1134 , \1135 ,         \1136 , \1137 , \1138 , \1139 , \1140 , \1141 , \1142 , \1143 , \1144 , \1145 ,         \1146 , \1147 , \1148 , \1149 , \1150 , \1151 , \1152 , \1153 , \1154 , \1155 ,         \1156 , \1157 , \1158 , \1159 , \1160 , \1161 , \1162 , \1163 , \1164 , \1165 ,         \1166 , \1167 , \1168 , \1169 , \1170 , \1171 , \1172 , \1173 , \1174 , \1175 ,         \1176 , \1177 , \1178 , \1179 , \1180 , \1181 , \1182 , \1183 , \1184 , \1185 ,         \1186 , \1187 , \1188 , \1189 , \1190 , \1191 , \1192 , \1193 , \1194 , \1195 ,         \1196 , \1197 , \1198 , \1199 , \1200 , \1201 , \1202 , \1203 , \1204 , \1205 ,         \1206 , \1207 , \1208 , \1209 , \1210 , \1211 , \1212 , \1213 , \1214 , \1215 ,         \1216 , \1217 , \1218 , \1219 , \1220 , \1221 , \1222 , \1223 , \1224 , \1225 ,         \1226 , \1227 , \1228 , \1229 , \1230 , \1231 , \1232 , \1233 , \1234 , \1235 ,         \1236 , \1237 , \1238 , \1239 , \1240 , \1241 , \1242 , \1243 , \1244 , \1245 ,         \1246 , \1247 , \1248 , \1249 , \1250 , \1251 , \1252 , \1253 , \1254 , \1255 ,         \1256 , \1257 , \1258 , \1259 , \1260 , \1261 , \1262 , \1263 , \1264 , \1265 ,         \1266 , \1267 , \1268 , \1269 , \1270 , \1271 , \1272 , \1273 , \1274 , \1275 ,         \1276 , \1277 , \1278 , \1279 , \1280 , \1281 , \1282 , \1283 , \1284 , \1285 ,         \1286 , \1287 , \1288 , \1289 , \1290 , \1291 , \1292 , \1293 , \1294 , \1295 ,         \1296 , \1297 , \1298 , \1299 , \1300 , \1301 , \1302 , \1303 , \1304 , \1305 ,         \1306 , \1307 , \1308 , \1309 , \1310 , \1311 , \1312 , \1313 , \1314 , \1315 ,         \1316 , \1317 , \1318 , \1319 , \1320 , \1321 , \1322 , \1323 , \1324 , \1325 ,         \1326 , \1327 , \1328 , \1329 , \1330 , \1331 , \1332 , \1333 , \1334 , \1335 ,         \1336 , \1337 , \1338 , \1339 , \1340 , \1341 , \1342 , \1343 , \1344 , \1345 ,         \1346 , \1347 , \1348 , \1349 , \1350 , \1351 , \1352 , \1353 , \1354 , \1355 ,         \1356 , \1357 , \1358 , \1359 , \1360 , \1361 , \1362 , \1363 , \1364 , \1365 ,         \1366 , \1367 , \1368 , \1369 , \1370 , \1371 , \1372 , \1373 , \1374 , \1375 ,         \1376 , \1377 , \1378 , \1379 , \1380 , \1381 , \1382 , \1383 , \1384 , \1385 ,         \1386 , \1387 , \1388 , \1389 , \1390 , \1391 , \1392 , \1393 , \1394 , \1395 ,         \1396 , \1397 , \1398 , \1399 , \1400 , \1401 , \1402 , \1403 , \1404 , \1405 ,         \1406 , \1407 , \1408 , \1409 , \1410 , \1411 , \1412 , \1413 , \1414 , \1415 ,         \1416 , \1417 , \1418 , \1419 , \1420 , \1421 , \1422 , \1423 , \1424 , \1425 ,         \1426 , \1427 , \1428 , \1429 , \1430 , \1431 , \1432 , \1433 , \1434 , \1435 ,         \1436 , \1437 , \1438 , \1439 , \1440 , \1441 , \1442 , \1443 , \1444 , \1445 ,         \1446 , \1447 , \1448 , \1449 , \1450 , \1451 , \1452 , \1453 , \1454 , \1455 ,         \1456 , \1457 , \1458 , \1459 , \1460 , \1461 , \1462 , \1463 , \1464 , \1465 ,         \1466 , \1467 , \1468 , \1469 , \1470 , \1471 , \1472 , \1473 , \1474 , \1475 ,         \1476 , \1477 , \1478 , \1479 , \1480 , \1481 , \1482 , \1483 , \1484 , \1485 ,         \1486 , \1487 , \1488 , \1489 , \1490 , \1491 , \1492 , \1493 , \1494 , \1495 ,         \1496 , \1497 , \1498 , \1499 , \1500 , \1501 , \1502 , \1503 , \1504 , \1505 ,         \1506 , \1507 , \1508 , \1509 , \1510 , \1511 , \1512 , \1513 , \1514 , \1515 ,         \1516 , \1517 , \1518 , \1519 , \1520 , \1521 , \1522 , \1523 , \1524 , \1525 ,         \1526 , \1527 , \1528 , \1529 , \1530 , \1531 , \1532 , \1533 , \1534 , \1535 ,         \1536 , \1537 , \1538 , \1539 , \1540 , \1541 , \1542 , \1543 , \1544 , \1545 ,         \1546 , \1547 , \1548 , \1549 , \1550 , \1551 , \1552 , \1553 , \1554 , \1555 ,         \1556 , \1557 , \1558 , \1559 , \1560 , \1561 , \1562 , \1563 , \1564 , \1565 ,         \1566 , \1567 , \1568 , \1569 , \1570 , \1571 , \1572 , \1573 , \1574 , \1575 ,         \1576 , \1577 , \1578 , \1579 , \1580 , \1581 , \1582 , \1583 , \1584 , \1585 ,         \1586 , \1587 , \1588 , \1589 , \1590 , \1591 , \1592 , \1593 , \1594 , \1595 ,         \1596 , \1597 , \1598 , \1599 , \1600 , \1601 , \1602 , \1603 , \1604 , \1605 ,         \1606 , \1607 , \1608 , \1609 , \1610 , \1611 , \1612 , \1613 , \1614 , \1615 ,         \1616 , \1617 , \1618 , \1619 , \1620 , \1621 , \1622 , \1623 , \1624 , \1625 ,         \1626 , \1627 , \1628 , \1629 , \1630 , \1631 , \1632 , \1633 , \1634 , \1635 ,         \1636 , \1637 , \1638 , \1639 , \1640 , \1641 , \1642 , \1643 , \1644 , \1645 ,         \1646 , \1647 , \1648 , \1649 , \1650 , \1651 , \1652 , \1653 , \1654 , \1655 ,         \1656 , \1657 , \1658 , \1659 , \1660 , \1661 , \1662 , \1663 , \1664 , \1665 ,         \1666 , \1667 , \1668 , \1669 , \1670 , \1671 , \1672 , \1673 , \1674 , \1675 ,         \1676 , \1677 , \1678 , \1679 , \1680 , \1681 , \1682 , \1683 , \1684 , \1685 ,         \1686 , \1687 , \1688 , \1689 , \1690 , \1691 , \1692 , \1693 , \1694 , \1695 ,         \1696 , \1697 , \1698 , \1699 , \1700 , \1701 , \1702 , \1703 , \1704 , \1705 ,         \1706 , \1707 , \1708 , \1709 , \1710 , \1711 , \1712 , \1713 , \1714 , \1715 ,         \1716 , \1717 , \1718 , \1719 , \1720 , \1721 , \1722 , \1723 , \1724 , \1725 ,         \1726 , \1727 , \1728 , \1729 , \1730 , \1731 , \1732 , \1733 , \1734 , \1735 ,         \1736 , \1737 , \1738 , \1739 , \1740 , \1741 , \1742 , \1743 , \1744 , \1745 ,         \1746 , \1747 , \1748 , \1749 , \1750 , \1751 , \1752 , \1753 , \1754 , \1755 ,         \1756 , \1757 , \1758 , \1759 , \1760 , \1761 , \1762 , \1763 , \1764 , \1765 ,         \1766 , \1767 , \1768 , \1769 , \1770 , \1771 , \1772 , \1773 , \1774 , \1775 ,         \1776 , \1777 , \1778 , \1779 , \1780 , \1781 , \1782 , \1783 , \1784 , \1785 ,         \1786 , \1787 , \1788 , \1789 , \1790 , \1791 , \1792 , \1793 , \1794 , \1795 ,         \1796 , \1797 , \1798 , \1799 , \1800 , \1801 , \1802 , \1803 , \1804 , \1805 ,         \1806 , \1807 , \1808 , \1809 , \1810 , \1811 , \1812 , \1813 , \1814 , \1815 ,         \1816 , \1817 , \1818 , \1819 , \1820 , \1821 , \1822 , \1823 , \1824 , \1825 ,         \1826 , \1827 , \1828 , \1829 , \1830 , \1831 , \1832 , \1833 , \1834 , \1835 ,         \1836 , \1837 , \1838 , \1839 , \1840 , \1841 , \1842 , \1843 , \1844 , \1845 ,         \1846 , \1847 , \1848 , \1849 , \1850 , \1851 , \1852 , \1853 , \1854 , \1855 ,         \1856 , \1857 , \1858 , \1859 , \1860 , \1861 , \1862 , \1863 , \1864 , \1865 ,         \1866 , \1867 , \1868 , \1869 , \1870 , \1871 , \1872 , \1873 , \1874 , \1875 ,         \1876 , \1877 , \1878 , \1879 , \1880 , \1881 , \1882 , \1883 , \1884 , \1885 ,         \1886 , \1887 , \1888 , \1889 , \1890 , \1891 , \1892 , \1893 , \1894 , \1895 ,         \1896 , \1897 , \1898 , \1899 , \1900 , \1901 , \1902 , \1903 , \1904 , \1905 ,         \1906 , \1907 , \1908 , \1909 , \1910 , \1911 , \1912 , \1913 , \1914 , \1915 ,         \1916 , \1917 , \1918 , \1919 , \1920 , \1921 , \1922 , \1923 , \1924 , \1925 ,         \1926 , \1927 , \1928 , \1929 , \1930 , \1931 , \1932 , \1933 , \1934 , \1935 ,         \1936 , \1937 , \1938 , \1939 , \1940 , \1941 , \1942 , \1943 , \1944 , \1945 ,         \1946 , \1947 , \1948 , \1949 , \1950 , \1951 , \1952 , \1953 , \1954 , \1955 ,         \1956 , \1957 , \1958 , \1959 , \1960 , \1961 , \1962 , \1963 , \1964 , \1965 ,         \1966 , \1967 , \1968 , \1969 , \1970 , \1971 , \1972 , \1973 , \1974 , \1975 ,         \1976 , \1977 , \1978 , \1979 , \1980 , \1981 , \1982 , \1983 , \1984 , \1985 ,         \1986 , \1987 , \1988 , \1989 , \1990 , \1991 , \1992 , \1993 , \1994 , \1995 ,         \1996 , \1997 , \1998 , \1999 , \2000 , \2001 , \2002 , \2003 , \2004 , \2005 ,         \2006 , \2007 , \2008 , \2009 , \2010 , \2011 , \2012 , \2013 , \2014 , \2015 ,         \2016 , \2017 , \2018 , \2019 , \2020 , \2021 , \2022 , \2023 , \2024 , \2025 ,         \2026 , \2027 , \2028 , \2029 , \2030 , \2031 , \2032 , \2033 , \2034 , \2035 ,         \2036 , \2037 , \2038 , \2039 , \2040 , \2041 , \2042 , \2043 , \2044 , \2045 ,         \2046 , \2047 , \2048 , \2049 , \2050 , \2051 , \2052 , \2053 , \2054 , \2055 ,         \2056 , \2057 , \2058 , \2059 , \2060 , \2061 , \2062 , \2063 , \2064 , \2065 ,         \2066 , \2067 , \2068 , \2069 , \2070 , \2071 , \2072 , \2073 , \2074 , \2075 ,         \2076 , \2077 , \2078 , \2079 , \2080 , \2081 , \2082 , \2083 , \2084 , \2085 ,         \2086 , \2087 , \2088 , \2089 , \2090 , \2091 , \2092 , \2093 , \2094 , \2095 ,         \2096 , \2097 , \2098 , \2099 , \2100 , \2101 , \2102 , \2103 , \2104 , \2105 ,         \2106 , \2107 , \2108 , \2109 , \2110 , \2111 , \2112 , \2113 , \2114 , \2115 ,         \2116 , \2117 , \2118 , \2119 , \2120 , \2121 , \2122 , \2123 , \2124 , \2125 ,         \2126 , \2127 , \2128 , \2129 , \2130 , \2131 , \2132 , \2133 , \2134 , \2135 ,         \2136 , \2137 , \2138 , \2139 , \2140 , \2141 , \2142 , \2143 , \2144 , \2145 ,         \2146 , \2147 , \2148 , \2149 , \2150 , \2151 , \2152 , \2153 , \2154 , \2155 ,         \2156 , \2157 , \2158 , \2159 , \2160 , \2161 , \2162 , \2163 , \2164 , \2165 ,         \2166 , \2167 , \2168 , \2169 , \2170 , \2171 , \2172 , \2173 , \2174 , \2175 ,         \2176 , \2177 , \2178 , \2179 , \2180 , \2181 , \2182 , \2183 , \2184 , \2185 ,         \2186 , \2187 , \2188 , \2189 , \2190 , \2191 , \2192 , \2193 , \2194 , \2195 ,         \2196 , \2197 , \2198 , \2199 , \2200 , \2201 , \2202 , \2203 , \2204 , \2205 ,         \2206 , \2207 , \2208 , \2209 , \2210 , \2211 , \2212 , \2213 , \2214 , \2215 ,         \2216 , \2217 , \2218 , \2219 , \2220 , \2221 , \2222 , \2223 , \2224 , \2225 ,         \2226 , \2227 , \2228 , \2229 , \2230 , \2231 , \2232 , \2233 , \2234 , \2235 ,         \2236 , \2237 , \2238 , \2239 , \2240 , \2241 , \2242 , \2243 , \2244 , \2245 ,         \2246 , \2247 , \2248 , \2249 , \2250 , \2251 , \2252 , \2253 , \2254 , \2255 ,         \2256 , \2257 , \2258 , \2259 , \2260 , \2261 , \2262 , \2263 , \2264 , \2265 ,         \2266 , \2267 , \2268 , \2269 , \2270 , \2271 , \2272 , \2273 , \2274 , \2275 ,         \2276 , \2277 , \2278 , \2279 , \2280 , \2281 , \2282 , \2283 , \2284 , \2285 ,         \2286 , \2287 , \2288 , \2289 , \2290 , \2291 , \2292 , \2293 , \2294 , \2295 ,         \2296 , \2297 , \2298 , \2299 , \2300 , \2301 , \2302 , \2303 , \2304 , \2305 ,         \2306 , \2307 , \2308 , \2309 , \2310 , \2311 , \2312 , \2313 , \2314 , \2315 ,         \2316 , \2317 , \2318 , \2319 , \2320 , \2321 , \2322 , \2323 , \2324 , \2325 ,         \2326 , \2327 , \2328 , \2329 , \2330 , \2331 , \2332 , \2333 , \2334 , \2335 ,         \2336 , \2337 , \2338 , \2339 , \2340 , \2341 , \2342 , \2343 , \2344 , \2345 ,         \2346 , \2347 , \2348 , \2349 , \2350 , \2351 , \2352 , \2353 , \2354 , \2355 ,         \2356 , \2357 , \2358 , \2359 , \2360 , \2361 , \2362 , \2363 , \2364 , \2365 ,         \2366 , \2367 , \2368 , \2369 , \2370 , \2371 , \2372 , \2373 , \2374 , \2375 ,         \2376 , \2377 , \2378 , \2379 , \2380 , \2381 , \2382 , \2383 , \2384 , \2385 ,         \2386 , \2387 , \2388 , \2389 , \2390 , \2391 , \2392 , \2393 , \2394 , \2395 ,         \2396 , \2397 , \2398 , \2399 , \2400 , \2401 , \2402 , \2403 , \2404 , \2405 ,         \2406 , \2407 , \2408 , \2409 , \2410 , \2411 , \2412 , \2413 , \2414 , \2415 ,         \2416 , \2417 , \2418 , \2419 , \2420 , \2421 , \2422 , \2423 , \2424 , \2425 ,         \2426 , \2427 , \2428 , \2429 , \2430 , \2431 , \2432 , \2433 , \2434 , \2435 ,         \2436 , \2437 , \2438 , \2439 , \2440 , \2441 , \2442 , \2443 , \2444 , \2445 ,         \2446 , \2447 , \2448 , \2449 , \2450 , \2451 , \2452 , \2453 , \2454 , \2455 ,         \2456 , \2457 , \2458 , \2459 , \2460 , \2461 , \2462 , \2463 , \2464 , \2465 ,         \2466 , \2467 , \2468 , \2469 , \2470 , \2471 , \2472 , \2473 , \2474 , \2475 ,         \2476 , \2477 , \2478 , \2479 , \2480 , \2481 , \2482 , \2483 , \2484 , \2485 ,         \2486 , \2487 , \2488 , \2489 , \2490 , \2491 , \2492 , \2493 , \2494 , \2495 ,         \2496 , \2497 , \2498 , \2499 , \2500 , \2501 , \2502 , \2503 , \2504 , \2505 ,         \2506 , \2507 , \2508 , \2509 , \2510 , \2511 , \2512 , \2513 , \2514 , \2515 ,         \2516 , \2517 , \2518 , \2519 , \2520 , \2521 , \2522 , \2523 , \2524 , \2525 ,         \2526 , \2527 , \2528 , \2529 , \2530 , \2531 , \2532 , \2533 , \2534 , \2535 ,         \2536 , \2537 , \2538 , \2539 , \2540 , \2541 , \2542 , \2543 , \2544 , \2545 ,         \2546 , \2547 , \2548 , \2549 , \2550 , \2551 , \2552 , \2553 , \2554 , \2555 ,         \2556 , \2557 , \2558 , \2559 , \2560 , \2561 , \2562 , \2563 , \2564 , \2565 ,         \2566 , \2567 , \2568 , \2569 , \2570 , \2571 , \2572 , \2573 , \2574 , \2575 ,         \2576 , \2577 , \2578 , \2579 , \2580 , \2581 , \2582 , \2583 , \2584 , \2585 ,         \2586 , \2587 , \2588 , \2589 , \2590 , \2591 , \2592 , \2593 , \2594 , \2595 ,         \2596 , \2597 , \2598 , \2599 , \2600 , \2601 , \2602 , \2603 , \2604 , \2605 ,         \2606 , \2607 , \2608 , \2609 , \2610 , \2611 , \2612 , \2613 , \2614 , \2615 ,         \2616 , \2617 , \2618 , \2619 , \2620 , \2621 , \2622 , \2623 , \2624 , \2625 ,         \2626 , \2627 , \2628 , \2629 , \2630 , \2631 , \2632 , \2633 , \2634 , \2635 ,         \2636 , \2637 , \2638 , \2639 , \2640 , \2641 , \2642 , \2643 , \2644 , \2645 ,         \2646 , \2647 , \2648 , \2649 , \2650 , \2651 , \2652 , \2653 , \2654 , \2655 ,         \2656 , \2657 , \2658 , \2659 , \2660 , \2661 , \2662 , \2663 , \2664 , \2665 ,         \2666 , \2667 , \2668 , \2669 , \2670 , \2671 , \2672 , \2673 , \2674 , \2675 ,         \2676 , \2677 , \2678 , \2679 , \2680 , \2681 , \2682 , \2683 , \2684 , \2685 ,         \2686 , \2687 , \2688 , \2689 , \2690 , \2691 , \2692 , \2693 , \2694 , \2695 ,         \2696 , \2697 , \2698 , \2699 , \2700 , \2701 , \2702 , \2703 , \2704 , \2705 ,         \2706 , \2707 , \2708 , \2709 , \2710 , \2711 , \2712 , \2713 , \2714 , \2715 ,         \2716 , \2717 , \2718 , \2719 , \2720 , \2721 , \2722 , \2723 , \2724 , \2725 ,         \2726 , \2727 , \2728 , \2729 , \2730 , \2731 , \2732 , \2733 , \2734 , \2735 ,         \2736 , \2737 , \2738 , \2739 , \2740 , \2741 , \2742 , \2743 , \2744 , \2745 ,         \2746 , \2747 , \2748 , \2749 , \2750 , \2751 , \2752 , \2753 , \2754 , \2755 ,         \2756 , \2757 , \2758 , \2759 , \2760 , \2761 , \2762 , \2763 , \2764 , \2765 ,         \2766 , \2767 , \2768 , \2769 , \2770 , \2771 , \2772 , \2773 , \2774 , \2775 ,         \2776 , \2777 , \2778 , \2779 , \2780 , \2781 , \2782 , \2783 , \2784 , \2785 ,         \2786 , \2787 , \2788 , \2789 , \2790 , \2791 , \2792 , \2793 , \2794 , \2795 ,         \2796 , \2797 , \2798 , \2799 , \2800 , \2801 , \2802 , \2803 , \2804 , \2805 ,         \2806 , \2807 , \2808 , \2809 , \2810 , \2811 , \2812 , \2813 , \2814 , \2815 ,         \2816 , \2817 , \2818 , \2819 , \2820 , \2821 , \2822 , \2823 , \2824 , \2825 ,         \2826 , \2827 , \2828 , \2829 , \2830 , \2831 , \2832 , \2833 , \2834 , \2835 ,         \2836 , \2837 , \2838 , \2839 , \2840 , \2841 , \2842 , \2843 , \2844 , \2845 ,         \2846 , \2847 , \2848 , \2849 , \2850 , \2851 , \2852 , \2853 , \2854 , \2855 ,         \2856 , \2857 , \2858 , \2859 , \2860 , \2861 , \2862 , \2863 , \2864 , \2865 ,         \2866 , \2867 , \2868 , \2869 , \2870 , \2871 , \2872 , \2873 , \2874 , \2875 ,         \2876 , \2877 , \2878 , \2879 , \2880 , \2881 , \2882 , \2883 , \2884 , \2885 ,         \2886 , \2887 , \2888 , \2889 , \2890 , \2891 , \2892 , \2893 , \2894 , \2895 ,         \2896 , \2897 , \2898 , \2899 , \2900 , \2901 , \2902 , \2903 , \2904 , \2905 ,         \2906 , \2907 , \2908 , \2909 , \2910 , \2911 , \2912 , \2913 , \2914 , \2915 ,         \2916 , \2917 , \2918 , \2919 , \2920 , \2921 , \2922 , \2923 , \2924 , \2925 ,         \2926 , \2927 , \2928 , \2929 , \2930 , \2931 , \2932 , \2933 , \2934 , \2935 ,         \2936 , \2937 , \2938 , \2939 , \2940 , \2941 , \2942 , \2943 , \2944 , \2945 ,         \2946 , \2947 , \2948 , \2949 , \2950 , \2951 , \2952 , \2953 , \2954 , \2955 ,         \2956 , \2957 , \2958 , \2959 , \2960 , \2961 , \2962 , \2963 , \2964 , \2965 ,         \2966 , \2967 , \2968 , \2969 , \2970 , \2971 , \2972 , \2973 , \2974 , \2975 ,         \2976 , \2977 , \2978 , \2979 , \2980 , \2981 , \2982 , \2983 , \2984 , \2985 ,         \2986 , \2987 , \2988 , \2989 , \2990 , \2991 , \2992 , \2993 , \2994 , \2995 ,         \2996 , \2997 , \2998 , \2999 , \3000 , \3001 , \3002 , \3003 , \3004 , \3005 ,         \3006 , \3007 , \3008 , \3009 , \3010 , \3011 , \3012 , \3013 , \3014 , \3015 ,         \3016 , \3017 , \3018 , \3019 , \3020 , \3021 , \3022 , \3023 , \3024 , \3025 ,         \3026 , \3027 , \3028 , \3029 , \3030 , \3031 , \3032 , \3033 , \3034 , \3035 ,         \3036 , \3037 , \3038 , \3039 , \3040 , \3041 , \3042 , \3043 , \3044 , \3045 ,         \3046 , \3047 , \3048 , \3049 , \3050 , \3051 , \3052 , \3053 , \3054 , \3055 ,         \3056 , \3057 , \3058 , \3059 , \3060 , \3061 , \3062 , \3063 , \3064 , \3065 ,         \3066 , \3067 , \3068 , \3069 , \3070 , \3071 , \3072 , \3073 , \3074 , \3075 ,         \3076 , \3077 , \3078 , \3079 , \3080 , \3081 , \3082 , \3083 , \3084 , \3085 ,         \3086 , \3087 , \3088 , \3089 , \3090 , \3091 , \3092 , \3093 , \3094 , \3095 ,         \3096 , \3097 , \3098 , \3099 , \3100 , \3101 , \3102 , \3103 , \3104 , \3105 ,         \3106 , \3107 , \3108 , \3109 , \3110 , \3111 , \3112 , \3113 , \3114 , \3115 ,         \3116 , \3117 , \3118 , \3119 , \3120 , \3121 , \3122 , \3123 , \3124 , \3125 ,         \3126 , \3127 , \3128 , \3129 , \3130 , \3131 , \3132 , \3133 , \3134 , \3135 ,         \3136 , \3137 , \3138 , \3139 , \3140 , \3141 , \3142 , \3143 , \3144 , \3145 ,         \3146 , \3147 , \3148 , \3149 , \3150 , \3151 , \3152 , \3153 , \3154 , \3155 ,         \3156 , \3157 , \3158 , \3159 , \3160 , \3161 , \3162 , \3163 , \3164 , \3165 ,         \3166 , \3167 , \3168 , \3169 , \3170 , \3171 , \3172 , \3173 , \3174 , \3175 ,         \3176 , \3177 , \3178 , \3179 , \3180 , \3181 , \3182 , \3183 , \3184 , \3185 ,         \3186 , \3187 , \3188 , \3189 , \3190 , \3191 , \3192 , \3193 , \3194 , \3195 ,         \3196 , \3197 , \3198 , \3199 , \3200 , \3201 , \3202 , \3203 , \3204 , \3205 ,         \3206 , \3207 , \3208 , \3209 , \3210 , \3211 , \3212 , \3213 , \3214 , \3215 ,         \3216 , \3217 , \3218 , \3219 , \3220 , \3221 , \3222 , \3223 , \3224 , \3225 ,         \3226 , \3227 , \3228 , \3229 , \3230 , \3231 , \3232 , \3233 , \3234 , \3235 ,         \3236 , \3237 , \3238 , \3239 , \3240 , \3241 , \3242 , \3243 , \3244 , \3245 ,         \3246 , \3247 , \3248 , \3249 , \3250 , \3251 , \3252 , \3253 , \3254 , \3255 ,         \3256 , \3257 , \3258 , \3259 , \3260 , \3261 , \3262 , \3263 , \3264 , \3265 ,         \3266 , \3267 , \3268 , \3269 , \3270 , \3271 , \3272 , \3273 , \3274 , \3275 ,         \3276 , \3277 , \3278 , \3279 , \3280 , \3281 , \3282 , \3283 , \3284 , \3285 ,         \3286 , \3287 , \3288 , \3289 , \3290 , \3291 , \3292 , \3293 , \3294 , \3295 ,         \3296 , \3297 , \3298 , \3299 , \3300 , \3301 , \3302 , \3303 , \3304 , \3305 ,         \3306 , \3307 , \3308 , \3309 , \3310 , \3311 , \3312 , \3313 , \3314 , \3315 ,         \3316 , \3317 , \3318 , \3319 , \3320 , \3321 , \3322 , \3323 , \3324 , \3325 ,         \3326 , \3327 , \3328 , \3329 , \3330 , \3331 , \3332 , \3333 , \3334 , \3335 ,         \3336 , \3337 , \3338 , \3339 , \3340 , \3341 , \3342 , \3343 , \3344 , \3345 ,         \3346 , \3347 , \3348 , \3349 , \3350 , \3351 , \3352 , \3353 , \3354 , \3355 ,         \3356 , \3357 , \3358 , \3359 , \3360 , \3361 , \3362 , \3363 , \3364 , \3365 ,         \3366 , \3367 , \3368 , \3369 , \3370 , \3371 , \3372 , \3373 , \3374 , \3375 ,         \3376 , \3377 , \3378 , \3379 , \3380 , \3381 , \3382 , \3383 , \3384 , \3385 ,         \3386 , \3387 , \3388 , \3389 , \3390 , \3391 , \3392 , \3393 , \3394 , \3395 ,         \3396 , \3397 , \3398 , \3399 , \3400 , \3401 , \3402 , \3403 , \3404 , \3405 ,         \3406 , \3407 , \3408 , \3409 , \3410 , \3411 , \3412 , \3413 , \3414 , \3415 ,         \3416 , \3417 , \3418 , \3419 , \3420 , \3421 , \3422 , \3423 , \3424 , \3425 ,         \3426 , \3427 , \3428 , \3429 , \3430 , \3431 , \3432 , \3433 , \3434 , \3435 ,         \3436 , \3437 , \3438 , \3439 , \3440 , \3441 , \3442 , \3443 , \3444 , \3445 ,         \3446 , \3447 , \3448 , \3449 , \3450 , \3451 , \3452 , \3453 , \3454 , \3455 ,         \3456 , \3457 , \3458 , \3459 , \3460 , \3461 , \3462 , \3463 , \3464 , \3465 ,         \3466 , \3467 , \3468 , \3469 , \3470 , \3471 , \3472 , \3473 , \3474 , \3475 ,         \3476 , \3477 , \3478 , \3479 , \3480 , \3481 , \3482 , \3483 , \3484 , \3485 ,         \3486 , \3487 , \3488 , \3489 , \3490 , \3491 , \3492 , \3493 , \3494 , \3495 ,         \3496 , \3497 , \3498 , \3499 , \3500 , \3501 , \3502 , \3503 , \3504 , \3505 ,         \3506 , \3507 , \3508 , \3509 , \3510 , \3511 , \3512 , \3513 , \3514 , \3515 ,         \3516 , \3517 , \3518 , \3519 , \3520 , \3521 , \3522 , \3523 , \3524 , \3525 ,         \3526 , \3527 , \3528 , \3529 , \3530 , \3531 , \3532 , \3533 , \3534 , \3535 ,         \3536 , \3537 , \3538 , \3539 , \3540 , \3541 , \3542 , \3543 , \3544 , \3545 ,         \3546 , \3547 , \3548 , \3549 , \3550 , \3551 , \3552 , \3553 , \3554 , \3555 ,         \3556 , \3557 , \3558 , \3559 , \3560 , \3561 , \3562 , \3563 , \3564 , \3565 ,         \3566 , \3567 , \3568 , \3569 , \3570 , \3571 , \3572 , \3573 , \3574 , \3575 ,         \3576 , \3577 , \3578 , \3579 , \3580 , \3581 , \3582 , \3583 , \3584 , \3585 ,         \3586 , \3587 , \3588 , \3589 , \3590 , \3591 , \3592 , \3593 , \3594 , \3595 ,         \3596 , \3597 , \3598 , \3599 , \3600 , \3601 , \3602 , \3603 , \3604 , \3605 ,         \3606 , \3607 , \3608 , \3609 , \3610 , \3611 , \3612 , \3613 , \3614 , \3615 ,         \3616 , \3617 , \3618 , \3619 , \3620 , \3621 , \3622 , \3623 , \3624 , \3625 ,         \3626 , \3627 , \3628 , \3629 , \3630 , \3631 , \3632 , \3633 , \3634 , \3635 ,         \3636 , \3637 , \3638 , \3639 , \3640 , \3641 , \3642 , \3643 , \3644 , \3645 ,         \3646 , \3647 , \3648 , \3649 , \3650 , \3651 , \3652 , \3653 , \3654 , \3655 ,         \3656 , \3657 , \3658 , \3659 , \3660 , \3661 , \3662 , \3663 , \3664 , \3665 ,         \3666 , \3667 , \3668 , \3669 , \3670 , \3671 , \3672 , \3673 , \3674 , \3675 ,         \3676 , \3677 , \3678 , \3679 , \3680 , \3681 , \3682 , \3683 , \3684 , \3685 ,         \3686 , \3687 , \3688 , \3689 , \3690 , \3691 , \3692 , \3693 , \3694 , \3695 ,         \3696 , \3697 , \3698 , \3699 , \3700 , \3701 , \3702 , \3703 , \3704 , \3705 ,         \3706 , \3707 , \3708 , \3709 , \3710 , \3711 , \3712 , \3713 , \3714 , \3715 ,         \3716 , \3717 , \3718 , \3719 , \3720 , \3721 , \3722 , \3723 , \3724 , \3725 ,         \3726 , \3727 , \3728 , \3729 , \3730 , \3731 , \3732 , \3733 , \3734 , \3735 ,         \3736 , \3737 , \3738 , \3739 , \3740 , \3741 , \3742 , \3743 , \3744 , \3745 ,         \3746 , \3747 , \3748 , \3749 , \3750 , \3751 , \3752 , \3753 , \3754 , \3755 ,         \3756 , \3757 , \3758 , \3759 , \3760 , \3761 , \3762 , \3763 , \3764 , \3765 ,         \3766 , \3767 , \3768 , \3769 , \3770 , \3771 , \3772 , \3773 , \3774 , \3775 ,         \3776 , \3777 , \3778 , \3779 , \3780 , \3781 , \3782 , \3783 , \3784 , \3785 ,         \3786 , \3787 , \3788 , \3789 , \3790 , \3791 , \3792 , \3793 , \3794 , \3795 ,         \3796 , \3797 , \3798 , \3799 , \3800 , \3801 , \3802 , \3803 , \3804 , \3805 ,         \3806 , \3807 , \3808 , \3809 , \3810 , \3811 , \3812 , \3813 , \3814 , \3815 ,         \3816 , \3817 , \3818 , \3819 , \3820 , \3821 , \3822 , \3823 , \3824 , \3825 ,         \3826 , \3827 , \3828 , \3829 , \3830 , \3831 , \3832 , \3833 , \3834 , \3835 ,         \3836 , \3837 , \3838 , \3839 , \3840 , \3841 , \3842 , \3843 , \3844 , \3845 ,         \3846 , \3847 , \3848 , \3849 , \3850 , \3851 , \3852 , \3853 , \3854 , \3855 ,         \3856 , \3857 , \3858 , \3859 , \3860 , \3861 , \3862 , \3863 , \3864 , \3865 ,         \3866 , \3867 , \3868 , \3869 , \3870 , \3871 , \3872 , \3873 , \3874 , \3875 ,         \3876 , \3877 , \3878 , \3879 , \3880 , \3881 , \3882 , \3883 , \3884 , \3885 ,         \3886 , \3887 , \3888 , \3889 , \3890 , \3891 , \3892 , \3893 , \3894 , \3895 ,         \3896 , \3897 , \3898 , \3899 , \3900 , \3901 , \3902 , \3903 , \3904 , \3905 ,         \3906 , \3907 , \3908 , \3909 , \3910 , \3911 , \3912 , \3913 , \3914 , \3915 ,         \3916 , \3917 , \3918 , \3919 , \3920 , \3921 , \3922 , \3923 , \3924 , \3925 ,         \3926 , \3927 , \3928 , \3929 , \3930 , \3931 , \3932 , \3933 , \3934 , \3935 ,         \3936 , \3937 , \3938 , \3939 , \3940 , \3941 , \3942 , \3943 , \3944 , \3945 ,         \3946 , \3947 , \3948 , \3949 , \3950 , \3951 , \3952 , \3953 , \3954 , \3955 ,         \3956 , \3957 , \3958 , \3959 , \3960 , \3961 , \3962 , \3963 , \3964 , \3965 ,         \3966 , \3967 , \3968 , \3969 , \3970 , \3971 , \3972 , \3973 , \3974 , \3975 ,         \3976 , \3977 , \3978 , \3979 , \3980 , \3981 , \3982 , \3983 , \3984 , \3985 ,         \3986 , \3987 , \3988 , \3989 , \3990 , \3991 , \3992 , \3993 , \3994 , \3995 ,         \3996 , \3997 , \3998 , \3999 , \4000 , \4001 , \4002 , \4003 , \4004 , \4005 ,         \4006 , \4007 , \4008 , \4009 , \4010 , \4011 , \4012 , \4013 , \4014 , \4015 ,         \4016 , \4017 , \4018 , \4019 , \4020 , \4021 , \4022 , \4023 , \4024 , \4025 ,         \4026 , \4027 , \4028 , \4029 , \4030 , \4031 , \4032 , \4033 , \4034 , \4035 ,         \4036 , \4037 , \4038 , \4039 , \4040 , \4041 , \4042 , \4043 , \4044 , \4045 ,         \4046 , \4047 , \4048 , \4049 , \4050 , \4051 , \4052 , \4053 , \4054 , \4055 ,         \4056 , \4057 , \4058 , \4059 , \4060 , \4061 , \4062 , \4063 , \4064 , \4065 ,         \4066 , \4067 , \4068 , \4069 , \4070 , \4071 , \4072 , \4073 , \4074 , \4075 ,         \4076 , \4077 , \4078 , \4079 , \4080 , \4081 , \4082 , \4083 , \4084 , \4085 ,         \4086 , \4087 , \4088 , \4089 , \4090 , \4091 , \4092 , \4093 , \4094 , \4095 ,         \4096 , \4097 , \4098 , \4099 , \4100 , \4101 , \4102 , \4103 , \4104 , \4105 ,         \4106 , \4107 , \4108 , \4109 , \4110 , \4111 , \4112 , \4113 , \4114 , \4115 ,         \4116 , \4117 , \4118 , \4119 , \4120 , \4121 , \4122 , \4123 , \4124 , \4125 ,         \4126 , \4127 , \4128 , \4129 , \4130 , \4131 , \4132 , \4133 , \4134 , \4135 ,         \4136 , \4137 , \4138 , \4139 , \4140 , \4141 , \4142 , \4143 , \4144 , \4145 ,         \4146 , \4147 , \4148 , \4149 , \4150 , \4151 , \4152 , \4153 , \4154 , \4155 ,         \4156 , \4157 , \4158 , \4159 , \4160 , \4161 , \4162 , \4163 , \4164 , \4165 ,         \4166 , \4167 , \4168 , \4169 , \4170 , \4171 , \4172 , \4173 , \4174 , \4175 ,         \4176 , \4177 , \4178 , \4179 , \4180 , \4181 , \4182 , \4183 , \4184 , \4185 ,         \4186 , \4187 , \4188 , \4189 , \4190 , \4191 , \4192 , \4193 , \4194 , \4195 ,         \4196 , \4197 , \4198 , \4199 , \4200 , \4201 , \4202 , \4203 , \4204 , \4205 ,         \4206 , \4207 , \4208 , \4209 , \4210 , \4211 , \4212 , \4213 , \4214 , \4215 ,         \4216 , \4217 , \4218 , \4219 , \4220 , \4221 , \4222 , \4223 , \4224 , \4225 ,         \4226 , \4227 , \4228 , \4229 , \4230 , \4231 , \4232 , \4233 , \4234 , \4235 ,         \4236 , \4237 , \4238 , \4239 , \4240 , \4241 , \4242 , \4243 , \4244 , \4245 ,         \4246 , \4247 , \4248 , \4249 , \4250 , \4251 , \4252 , \4253 , \4254 , \4255 ,         \4256 , \4257 , \4258 , \4259 , \4260 , \4261 , \4262 , \4263 , \4264 , \4265 ,         \4266 , \4267 , \4268 , \4269 , \4270 , \4271 , \4272 , \4273 , \4274 , \4275 ,         \4276 , \4277 , \4278 , \4279 , \4280 , \4281 , \4282 , \4283 , \4284 , \4285 ,         \4286 , \4287 , \4288 , \4289 , \4290 , \4291 , \4292 , \4293 , \4294 , \4295 ,         \4296 , \4297 , \4298 , \4299 , \4300 , \4301 , \4302 , \4303 , \4304 , \4305 ,         \4306 , \4307 , \4308 , \4309 , \4310 , \4311 , \4312 , \4313 , \4314 , \4315 ,         \4316 , \4317 , \4318 , \4319 , \4320 , \4321 , \4322 , \4323 , \4324 , \4325 ,         \4326 , \4327 , \4328 , \4329 , \4330 , \4331 , \4332 , \4333 , \4334 , \4335 ,         \4336 , \4337 , \4338 , \4339 , \4340 , \4341 , \4342 , \4343 , \4344 , \4345 ,         \4346 , \4347 , \4348 , \4349 , \4350 , \4351 , \4352 , \4353 , \4354 , \4355 ,         \4356 , \4357 , \4358 , \4359 , \4360 , \4361 , \4362 , \4363 , \4364 , \4365 ,         \4366 , \4367 , \4368 , \4369 , \4370 , \4371 , \4372 , \4373 , \4374 , \4375 ,         \4376 , \4377 , \4378 , \4379 , \4380 , \4381 , \4382 , \4383 , \4384 , \4385 ,         \4386 , \4387 , \4388 , \4389 , \4390 , \4391 , \4392 , \4393 , \4394 , \4395 ,         \4396 , \4397 , \4398 , \4399 , \4400 , \4401 , \4402 , \4403 , \4404 , \4405 ,         \4406 , \4407 , \4408 , \4409 , \4410 , \4411 , \4412 , \4413 , \4414 , \4415 ,         \4416 , \4417 , \4418 , \4419 , \4420 , \4421 , \4422 , \4423 , \4424 , \4425 ,         \4426 , \4427 , \4428 , \4429 , \4430 , \4431 , \4432 , \4433 , \4434 , \4435 ,         \4436 , \4437 , \4438 , \4439 , \4440 , \4441 , \4442 , \4443 , \4444 , \4445 ,         \4446 , \4447 , \4448 , \4449 , \4450 , \4451 , \4452 , \4453 , \4454 , \4455 ,         \4456 , \4457 , \4458 , \4459 , \4460 , \4461 , \4462 , \4463 , \4464 , \4465 ,         \4466 , \4467 , \4468 , \4469 , \4470 , \4471 , \4472 , \4473 , \4474 , \4475 ,         \4476 , \4477 , \4478 , \4479 , \4480 , \4481 , \4482 , \4483 , \4484 , \4485 ,         \4486 , \4487 , \4488 , \4489 , \4490 , \4491 , \4492 , \4493 , \4494 , \4495 ,         \4496 , \4497 , \4498 , \4499 , \4500 , \4501 , \4502 , \4503 , \4504 , \4505 ,         \4506 , \4507 , \4508 , \4509 , \4510 , \4511 , \4512 , \4513 , \4514 , \4515 ,         \4516 , \4517 , \4518 , \4519 , \4520 , \4521 , \4522 , \4523 , \4524 , \4525 ,         \4526 , \4527 , \4528 , \4529 , \4530 , \4531 , \4532 , \4533 , \4534 , \4535 ,         \4536 , \4537 , \4538 , \4539 , \4540 , \4541 , \4542 , \4543 , \4544 , \4545 ,         \4546 , \4547 , \4548 , \4549 , \4550 , \4551 , \4552 , \4553 , \4554 , \4555 ,         \4556 , \4557 , \4558 , \4559 , \4560 , \4561 , \4562 , \4563 , \4564 , \4565 ,         \4566 , \4567 , \4568 , \4569 , \4570 , \4571 , \4572 , \4573 , \4574 , \4575 ,         \4576 , \4577 , \4578 , \4579 , \4580 , \4581 , \4582 , \4583 , \4584 , \4585 ,         \4586 , \4587 , \4588 , \4589 , \4590 , \4591 , \4592 , \4593 , \4594 , \4595 ,         \4596 , \4597 , \4598 , \4599 , \4600 , \4601 , \4602 , \4603 , \4604 , \4605 ,         \4606 , \4607 , \4608 , \4609 , \4610 , \4611 , \4612 , \4613 , \4614 , \4615 ,         \4616 , \4617 , \4618 , \4619 , \4620 , \4621 , \4622 , \4623 , \4624 , \4625 ,         \4626 , \4627 , \4628 , \4629 , \4630 , \4631 , \4632 , \4633 , \4634 , \4635 ,         \4636 , \4637 , \4638 , \4639 , \4640 , \4641 , \4642 , \4643 , \4644 , \4645 ,         \4646 , \4647 , \4648 , \4649 , \4650 , \4651 , \4652 , \4653 , \4654 , \4655 ,         \4656 , \4657 , \4658 , \4659 , \4660 , \4661 , \4662 , \4663 , \4664 , \4665 ,         \4666 , \4667 , \4668 , \4669 , \4670 , \4671 , \4672 , \4673 , \4674 , \4675 ,         \4676 , \4677 , \4678 , \4679 , \4680 , \4681 , \4682 , \4683 , \4684 , \4685 ,         \4686 , \4687 , \4688 , \4689 , \4690 , \4691 , \4692 , \4693 , \4694 , \4695 ,         \4696 , \4697 , \4698 , \4699 , \4700 , \4701 , \4702 , \4703 , \4704 , \4705 ,         \4706 , \4707 , \4708 , \4709 , \4710 , \4711 , \4712 , \4713 , \4714 , \4715 ,         \4716 , \4717 , \4718 , \4719 , \4720 , \4721 , \4722 , \4723 , \4724 , \4725 ,         \4726 , \4727 , \4728 , \4729 , \4730 , \4731 , \4732 , \4733 , \4734 , \4735 ,         \4736 , \4737 , \4738 , \4739 , \4740 , \4741 , \4742 , \4743 , \4744 , \4745 ,         \4746 , \4747 , \4748 , \4749 , \4750 , \4751 , \4752 , \4753 , \4754 , \4755 ,         \4756 , \4757 , \4758 , \4759 , \4760 , \4761 , \4762 , \4763 , \4764 , \4765 ,         \4766 , \4767 , \4768 , \4769 , \4770 , \4771 , \4772 , \4773 , \4774 , \4775 ,         \4776 , \4777 , \4778 , \4779 , \4780 , \4781 , \4782 , \4783 , \4784 , \4785 ,         \4786 , \4787 , \4788 , \4789 , \4790 , \4791 , \4792 , \4793 , \4794 , \4795 ,         \4796 , \4797 , \4798 , \4799 , \4800 , \4801 , \4802 , \4803 , \4804 , \4805 ,         \4806 , \4807 , \4808 , \4809 , \4810 , \4811 , \4812 , \4813 , \4814 , \4815 ,         \4816 , \4817 , \4818 , \4819 , \4820 , \4821 , \4822 , \4823 , \4824 , \4825 ,         \4826 , \4827 , \4828 , \4829 , \4830 , \4831 , \4832 , \4833 , \4834 , \4835 ,         \4836 , \4837 , \4838 , \4839 , \4840 , \4841 , \4842 , \4843 , \4844 , \4845 ,         \4846 , \4847 , \4848 , \4849 , \4850 , \4851 , \4852 , \4853 , \4854 , \4855 ,         \4856 , \4857 , \4858 , \4859 , \4860 , \4861 , \4862 , \4863 , \4864 , \4865 ,         \4866 , \4867 , \4868 , \4869 , \4870 , \4871 , \4872 , \4873 , \4874 , \4875 ,         \4876 , \4877 , \4878 , \4879 , \4880 , \4881 , \4882 , \4883 , \4884 , \4885 ,         \4886 , \4887 , \4888 , \4889 , \4890 , \4891 , \4892 , \4893 , \4894 , \4895 ,         \4896 , \4897 , \4898 , \4899 , \4900 , \4901 , \4902 , \4903 , \4904 , \4905 ,         \4906 , \4907 , \4908 , \4909 , \4910 , \4911 , \4912 , \4913 , \4914 , \4915 ,         \4916 , \4917 , \4918 , \4919 , \4920 , \4921 , \4922 , \4923 , \4924 , \4925 ,         \4926 , \4927 , \4928 , \4929 , \4930 , \4931 , \4932 , \4933 , \4934 , \4935 ,         \4936 , \4937 , \4938 , \4939 , \4940 , \4941 , \4942 , \4943 , \4944 , \4945 ,         \4946 , \4947 , \4948 , \4949 , \4950 , \4951 , \4952 , \4953 , \4954 , \4955 ,         \4956 , \4957 , \4958 , \4959 , \4960 , \4961 , \4962 , \4963 , \4964 , \4965 ,         \4966 , \4967 , \4968 , \4969 , \4970 , \4971 , \4972 , \4973 , \4974 , \4975 ,         \4976 , \4977 , \4978 , \4979 , \4980 , \4981 , \4982 , \4983 , \4984 , \4985 ,         \4986 , \4987 , \4988 , \4989 , \4990 , \4991 , \4992 , \4993 , \4994 , \4995 ,         \4996 , \4997 , \4998 , \4999 , \5000 , \5001 , \5002 , \5003 , \5004 , \5005 ,         \5006 , \5007 , \5008 , \5009 , \5010 , \5011 , \5012 , \5013 , \5014 , \5015 ,         \5016 , \5017 , \5018 , \5019 , \5020 , \5021 , \5022 , \5023 , \5024 , \5025 ,         \5026 , \5027 , \5028 , \5029 , \5030 , \5031 , \5032 , \5033 , \5034 , \5035 ,         \5036 , \5037 , \5038 , \5039 , \5040 , \5041 , \5042 , \5043 , \5044 , \5045 ,         \5046 , \5047 , \5048 , \5049 , \5050 , \5051 , \5052 , \5053 , \5054 , \5055 ,         \5056 , \5057 , \5058 , \5059 , \5060 , \5061 , \5062 , \5063 , \5064 , \5065 ,         \5066 , \5067 , \5068 , \5069 , \5070 , \5071 , \5072 , \5073 , \5074 , \5075 ,         \5076 , \5077 , \5078 , \5079 , \5080 , \5081 , \5082 , \5083 , \5084 , \5085 ,         \5086 , \5087 , \5088 , \5089 , \5090 , \5091 , \5092 , \5093 , \5094 , \5095 ,         \5096 , \5097 , \5098 , \5099 , \5100 , \5101 , \5102 , \5103 , \5104 , \5105 ,         \5106 , \5107 , \5108 , \5109 , \5110 , \5111 , \5112 , \5113 , \5114 , \5115 ,         \5116 , \5117 , \5118 , \5119 , \5120 , \5121 , \5122 , \5123 , \5124 , \5125 ,         \5126 , \5127 , \5128 , \5129 , \5130 , \5131 , \5132 , \5133 , \5134 , \5135 ,         \5136 , \5137 , \5138 , \5139 , \5140 , \5141 , \5142 , \5143 , \5144 , \5145 ,         \5146 , \5147 , \5148 , \5149 , \5150 , \5151 , \5152 , \5153 , \5154 , \5155 ,         \5156 , \5157 , \5158 , \5159 , \5160 , \5161 , \5162 , \5163 , \5164 , \5165 ,         \5166 , \5167 , \5168 , \5169 , \5170 , \5171 , \5172 , \5173 , \5174 , \5175 ,         \5176 , \5177 , \5178 , \5179 , \5180 , \5181 , \5182 , \5183 , \5184 , \5185 ,         \5186 , \5187 , \5188 , \5189 , \5190 , \5191 , \5192 , \5193 , \5194 , \5195 ,         \5196 , \5197 , \5198 , \5199 , \5200 , \5201 , \5202 , \5203 , \5204 , \5205 ,         \5206 , \5207 , \5208 , \5209 , \5210 , \5211 , \5212 , \5213 , \5214 , \5215 ,         \5216 , \5217 , \5218 , \5219 , \5220 , \5221 , \5222 , \5223 , \5224 , \5225 ,         \5226 , \5227 , \5228 , \5229 , \5230 , \5231 , \5232 , \5233 , \5234 , \5235 ,         \5236 , \5237 , \5238 , \5239 , \5240 , \5241 , \5242 , \5243 , \5244 , \5245 ,         \5246 , \5247 , \5248 , \5249 , \5250 , \5251 , \5252 , \5253 , \5254 , \5255 ,         \5256 , \5257 , \5258 , \5259 , \5260 , \5261 , \5262 , \5263 , \5264 , \5265 ,         \5266 , \5267 , \5268 , \5269 , \5270 , \5271 , \5272 , \5273 , \5274 , \5275 ,         \5276 , \5277 , \5278 , \5279 , \5280 , \5281 , \5282 , \5283 , \5284 , \5285 ,         \5286 , \5287 , \5288 , \5289 , \5290 , \5291 , \5292 , \5293 , \5294 , \5295 ,         \5296 , \5297 , \5298 , \5299 , \5300 , \5301 , \5302 , \5303 , \5304 , \5305 ,         \5306 , \5307 , \5308 , \5309 , \5310 , \5311 , \5312 , \5313 , \5314 , \5315 ,         \5316 , \5317 , \5318 , \5319 , \5320 , \5321 , \5322 , \5323 , \5324 , \5325 ,         \5326 , \5327 , \5328 , \5329 , \5330 , \5331 , \5332 , \5333 , \5334 , \5335 ,         \5336 , \5337 , \5338 , \5339 , \5340 , \5341 , \5342 , \5343 , \5344 , \5345 ,         \5346 , \5347 , \5348 , \5349 , \5350 , \5351 , \5352 , \5353 , \5354 , \5355 ,         \5356 , \5357 , \5358 , \5359 , \5360 , \5361 , \5362 , \5363 , \5364 , \5365 ,         \5366 , \5367 , \5368 , \5369 , \5370 , \5371 , \5372 , \5373 , \5374 , \5375 ,         \5376 , \5377 , \5378 , \5379 , \5380 , \5381 , \5382 , \5383 , \5384 , \5385 ,         \5386 , \5387 , \5388 , \5389 , \5390 , \5391 , \5392 , \5393 , \5394 , \5395 ,         \5396 , \5397 , \5398 , \5399 , \5400 , \5401 , \5402 , \5403 , \5404 , \5405 ,         \5406 , \5407 , \5408 , \5409 , \5410 , \5411 , \5412 , \5413 , \5414 , \5415 ,         \5416 , \5417 , \5418 , \5419 , \5420 , \5421 , \5422 , \5423 , \5424 , \5425 ,         \5426 , \5427 , \5428 , \5429 , \5430 , \5431 , \5432 , \5433 , \5434 , \5435 ,         \5436 , \5437 , \5438 , \5439 , \5440 , \5441 , \5442 , \5443 , \5444 , \5445 ,         \5446 , \5447 , \5448 , \5449 , \5450 , \5451 , \5452 , \5453 , \5454 , \5455 ,         \5456 , \5457 , \5458 , \5459 , \5460 , \5461 , \5462 , \5463 , \5464 , \5465 ,         \5466 , \5467 , \5468 , \5469 , \5470 , \5471 , \5472 , \5473 , \5474 , \5475 ,         \5476 , \5477 , \5478 , \5479 , \5480 , \5481 , \5482 , \5483 , \5484 , \5485 ,         \5486 , \5487 , \5488 , \5489 , \5490 , \5491 , \5492 , \5493 , \5494 , \5495 ,         \5496 , \5497 , \5498 , \5499 , \5500 , \5501 , \5502 , \5503 , \5504 , \5505 ,         \5506 , \5507 , \5508 , \5509 , \5510 , \5511 , \5512 , \5513 , \5514 , \5515 ,         \5516 , \5517 , \5518 , \5519 , \5520 , \5521 , \5522 , \5523 , \5524 , \5525 ,         \5526 , \5527 , \5528 , \5529 , \5530 , \5531 , \5532 , \5533 , \5534 , \5535 ,         \5536 , \5537 , \5538 , \5539 , \5540 , \5541 , \5542 , \5543 , \5544 , \5545 ,         \5546 , \5547 , \5548 , \5549 , \5550 , \5551 , \5552 , \5553 , \5554 , \5555 ,         \5556 , \5557 , \5558 , \5559 , \5560 , \5561 , \5562 , \5563 , \5564 , \5565 ,         \5566 , \5567 , \5568 , \5569 , \5570 , \5571 , \5572 , \5573 , \5574 , \5575 ,         \5576 , \5577 , \5578 , \5579 , \5580 , \5581 , \5582 , \5583 , \5584 , \5585 ,         \5586 , \5587 , \5588 , \5589 , \5590 , \5591 , \5592 , \5593 , \5594 , \5595 ,         \5596 , \5597 , \5598 , \5599 , \5600 , \5601 , \5602 , \5603 , \5604 , \5605 ,         \5606 , \5607 , \5608 , \5609 , \5610 , \5611 , \5612 , \5613 , \5614 , \5615 ,         \5616 , \5617 , \5618 , \5619 , \5620 , \5621 , \5622 , \5623 , \5624 , \5625 ,         \5626 , \5627 , \5628 , \5629 , \5630 , \5631 , \5632 , \5633 , \5634 , \5635 ,         \5636 , \5637 , \5638 , \5639 , \5640 , \5641 , \5642 , \5643 , \5644 , \5645 ,         \5646 , \5647 , \5648 , \5649 , \5650 , \5651 , \5652 , \5653 , \5654 , \5655 ,         \5656 , \5657 , \5658 , \5659 , \5660 , \5661 , \5662 , \5663 , \5664 , \5665 ,         \5666 , \5667 , \5668 , \5669 , \5670 , \5671 , \5672 , \5673 , \5674 , \5675 ,         \5676 , \5677 , \5678 , \5679 , \5680 , \5681 , \5682 , \5683 , \5684 , \5685 ,         \5686 , \5687 , \5688 , \5689 , \5690 , \5691 , \5692 , \5693 , \5694 , \5695 ,         \5696 , \5697 , \5698 , \5699 , \5700 , \5701 , \5702 , \5703 , \5704 , \5705 ,         \5706 , \5707 , \5708 , \5709 , \5710 , \5711 , \5712 , \5713 , \5714 , \5715 ,         \5716 , \5717 , \5718 , \5719 , \5720 , \5721 , \5722 , \5723 , \5724 , \5725 ,         \5726 , \5727 , \5728 , \5729 , \5730 , \5731 , \5732 , \5733 , \5734 , \5735 ,         \5736 , \5737 , \5738 , \5739 , \5740 , \5741 , \5742 , \5743 , \5744 , \5745 ,         \5746 , \5747 , \5748 , \5749 , \5750 , \5751 , \5752 , \5753 , \5754 , \5755 ,         \5756 , \5757 , \5758 , \5759 , \5760 , \5761 , \5762 , \5763 , \5764 , \5765 ,         \5766 , \5767 , \5768 , \5769 , \5770 , \5771 , \5772 , \5773 , \5774 , \5775 ,         \5776 , \5777 , \5778 , \5779 , \5780 , \5781 , \5782 , \5783 , \5784 , \5785 ,         \5786 , \5787 , \5788 , \5789 , \5790 , \5791 , \5792 , \5793 , \5794 , \5795 ,         \5796 , \5797 , \5798 , \5799 , \5800 , \5801 , \5802 , \5803 , \5804 , \5805 ,         \5806 , \5807 , \5808 , \5809 , \5810 , \5811 , \5812 , \5813 , \5814 , \5815 ,         \5816 , \5817 , \5818 , \5819 , \5820 , \5821 , \5822 , \5823 , \5824 , \5825 ,         \5826 , \5827 , \5828 , \5829 , \5830 , \5831 , \5832 , \5833 , \5834 , \5835 ,         \5836 , \5837 , \5838 , \5839 , \5840 , \5841 , \5842 , \5843 , \5844 , \5845 ,         \5846 , \5847 , \5848 , \5849 , \5850 , \5851 , \5852 , \5853 , \5854 , \5855 ,         \5856 , \5857 , \5858 , \5859 , \5860 , \5861 , \5862 , \5863 , \5864 , \5865 ,         \5866 , \5867 , \5868 , \5869 , \5870 , \5871 , \5872 , \5873 , \5874 , \5875 ,         \5876 , \5877 , \5878 , \5879 , \5880 , \5881 , \5882 , \5883 , \5884 , \5885 ,         \5886 , \5887 , \5888 , \5889 , \5890 , \5891 , \5892 , \5893 , \5894 , \5895 ,         \5896 , \5897 , \5898 , \5899 , \5900 , \5901 , \5902 , \5903 , \5904 , \5905 ,         \5906 , \5907 , \5908 , \5909 , \5910 , \5911 , \5912 , \5913 , \5914 , \5915 ,         \5916 , \5917 , \5918 , \5919 , \5920 , \5921 , \5922 , \5923 , \5924 , \5925 ,         \5926 , \5927 , \5928 , \5929 , \5930 , \5931 , \5932 , \5933 , \5934 , \5935 ,         \5936 , \5937 , \5938 , \5939 , \5940 , \5941 , \5942 , \5943 , \5944 , \5945 ,         \5946 , \5947 , \5948 , \5949 , \5950 , \5951 , \5952 , \5953 , \5954 , \5955 ,         \5956 , \5957 , \5958 , \5959 , \5960 , \5961 , \5962 , \5963 , \5964 , \5965 ,         \5966 , \5967 , \5968 , \5969 , \5970 , \5971 , \5972 , \5973 , \5974 , \5975 ,         \5976 , \5977 , \5978 , \5979 , \5980 , \5981 , \5982 , \5983 , \5984 , \5985 ,         \5986 , \5987 , \5988 , \5989 , \5990 , \5991 , \5992 , \5993 , \5994 , \5995 ,         \5996 , \5997 , \5998 , \5999 , \6000 , \6001 , \6002 , \6003 , \6004 , \6005 ,         \6006 , \6007 , \6008 , \6009 , \6010 , \6011 , \6012 , \6013 , \6014 , \6015 ,         \6016 , \6017 , \6018 , \6019 , \6020 , \6021 , \6022 , \6023 , \6024 , \6025 ,         \6026 , \6027 , \6028 , \6029 , \6030 , \6031 , \6032 , \6033 , \6034 , \6035 ,         \6036 , \6037 , \6038 , \6039 , \6040 , \6041 , \6042 , \6043 , \6044 , \6045 ,         \6046 , \6047 , \6048 , \6049 , \6050 , \6051 , \6052 , \6053 , \6054 , \6055 ,         \6056 , \6057 , \6058 , \6059 , \6060 , \6061 , \6062 , \6063 , \6064 , \6065 ,         \6066 , \6067 , \6068 , \6069 , \6070 , \6071 , \6072 , \6073 , \6074 , \6075 ,         \6076 , \6077 , \6078 , \6079 , \6080 , \6081 , \6082 , \6083 , \6084 , \6085 ,         \6086 , \6087 , \6088 , \6089 , \6090 , \6091 , \6092 , \6093 , \6094 , \6095 ,         \6096 , \6097 , \6098 , \6099 , \6100 , \6101 , \6102 , \6103 , \6104 , \6105 ,         \6106 , \6107 , \6108 , \6109 , \6110 , \6111 , \6112 , \6113 , \6114 , \6115 ,         \6116 , \6117 , \6118 , \6119 , \6120 , \6121 , \6122 , \6123 , \6124 , \6125 ,         \6126 , \6127 , \6128 , \6129 , \6130 , \6131 , \6132 , \6133 , \6134 , \6135 ,         \6136 , \6137 , \6138 , \6139 , \6140 , \6141 , \6142 , \6143 , \6144 , \6145 ,         \6146 , \6147 , \6148 , \6149 , \6150 , \6151 , \6152 , \6153 , \6154 , \6155 ,         \6156 , \6157 , \6158 , \6159 , \6160 , \6161 , \6162 , \6163 , \6164 , \6165 ,         \6166 , \6167 , \6168 , \6169 , \6170 , \6171 , \6172 , \6173 , \6174 , \6175 ,         \6176 , \6177 , \6178 , \6179 , \6180 , \6181 , \6182 , \6183 , \6184 , \6185 ,         \6186 , \6187 , \6188 , \6189 , \6190 , \6191 , \6192 , \6193 , \6194 , \6195 ,         \6196 , \6197 , \6198 , \6199 , \6200 , \6201 , \6202 , \6203 , \6204 , \6205 ,         \6206 , \6207 , \6208 , \6209 , \6210 , \6211 , \6212 , \6213 , \6214 , \6215 ,         \6216 , \6217 , \6218 , \6219 , \6220 , \6221 , \6222 , \6223 , \6224 , \6225 ,         \6226 , \6227 , \6228 , \6229 , \6230 , \6231 , \6232 , \6233 , \6234 , \6235 ,         \6236 , \6237 , \6238 , \6239 , \6240 , \6241 , \6242 , \6243 , \6244 , \6245 ,         \6246 , \6247 , \6248 , \6249 , \6250 , \6251 , \6252 , \6253 , \6254 , \6255 ,         \6256 , \6257 , \6258 , \6259 , \6260 , \6261 , \6262 , \6263 , \6264 , \6265 ,         \6266 , \6267 , \6268 , \6269 , \6270 , \6271 , \6272 , \6273 , \6274 , \6275 ,         \6276 , \6277 , \6278 , \6279 , \6280 , \6281 , \6282 , \6283 , \6284 , \6285 ,         \6286 , \6287 , \6288 , \6289 , \6290 , \6291 , \6292 , \6293 , \6294 , \6295 ,         \6296 , \6297 , \6298 , \6299 , \6300 , \6301 , \6302 , \6303 , \6304 , \6305 ,         \6306 , \6307 , \6308 , \6309 , \6310 , \6311 , \6312 , \6313 , \6314 , \6315 ,         \6316 , \6317 , \6318 , \6319 , \6320 , \6321 , \6322 , \6323 , \6324 , \6325 ,         \6326 , \6327 , \6328 , \6329 , \6330 , \6331 , \6332 , \6333 , \6334 , \6335 ,         \6336 , \6337 , \6338 , \6339 , \6340 , \6341 , \6342 , \6343 , \6344 , \6345 ,         \6346 , \6347 , \6348 , \6349 , \6350 , \6351 , \6352 , \6353 , \6354 , \6355 ,         \6356 , \6357 , \6358 , \6359 , \6360 , \6361 , \6362 , \6363 , \6364 , \6365 ,         \6366 , \6367 , \6368 , \6369 , \6370 , \6371 , \6372 , \6373 , \6374 , \6375 ,         \6376 , \6377 , \6378 , \6379 , \6380 , \6381 , \6382 , \6383 , \6384 , \6385 ,         \6386 , \6387 , \6388 , \6389 , \6390 , \6391 , \6392 , \6393 , \6394 , \6395 ,         \6396 , \6397 , \6398 , \6399 , \6400 , \6401 , \6402 , \6403 , \6404 , \6405 ,         \6406 , \6407 , \6408 , \6409 , \6410 , \6411 , \6412 , \6413 , \6414 , \6415 ,         \6416 , \6417 , \6418 , \6419 , \6420 , \6421 , \6422 , \6423 , \6424 , \6425 ,         \6426 , \6427 , \6428 , \6429 , \6430 , \6431 , \6432 , \6433 , \6434 , \6435 ,         \6436 , \6437 , \6438 , \6439 , \6440 , \6441 , \6442 , \6443 , \6444 , \6445 ,         \6446 , \6447 , \6448 , \6449 , \6450 , \6451 , \6452 , \6453 , \6454 , \6455 ,         \6456 , \6457 , \6458 , \6459 , \6460 , \6461 , \6462 , \6463 , \6464 , \6465 ,         \6466 , \6467 , \6468 , \6469 , \6470 , \6471 , \6472 , \6473 , \6474 , \6475 ,         \6476 , \6477 , \6478 , \6479 , \6480 , \6481 , \6482 , \6483 , \6484 , \6485 ,         \6486 , \6487 , \6488 , \6489 , \6490 , \6491 , \6492 , \6493 , \6494 , \6495 ,         \6496 , \6497 , \6498 , \6499 , \6500 , \6501 , \6502 , \6503 , \6504 , \6505 ,         \6506 , \6507 , \6508 , \6509 , \6510 , \6511 , \6512 , \6513 , \6514 , \6515 ,         \6516 , \6517 , \6518 , \6519 , \6520 , \6521 , \6522 , \6523 , \6524 , \6525 ,         \6526 , \6527 , \6528 , \6529 , \6530 , \6531 , \6532 , \6533 , \6534 , \6535 ,         \6536 , \6537 , \6538 , \6539 , \6540 , \6541 , \6542 , \6543 , \6544 , \6545 ,         \6546 , \6547 , \6548 , \6549 , \6550 , \6551 , \6552 , \6553 , \6554 , \6555 ,         \6556 , \6557 , \6558 , \6559 , \6560 , \6561 , \6562 , \6563 , \6564 , \6565 ,         \6566 , \6567 , \6568 , \6569 , \6570 , \6571 , \6572 , \6573 , \6574 , \6575 ,         \6576 , \6577 , \6578 , \6579 , \6580 , \6581 , \6582 , \6583 , \6584 , \6585 ,         \6586 , \6587 , \6588 , \6589 , \6590 , \6591 , \6592 , \6593 , \6594 , \6595 ,         \6596 , \6597 , \6598 , \6599 , \6600 , \6601 , \6602 , \6603 , \6604 , \6605 ,         \6606 , \6607 , \6608 , \6609 , \6610 , \6611 , \6612 , \6613 , \6614 , \6615 ,         \6616 , \6617 , \6618 , \6619 , \6620 , \6621 , \6622 , \6623 , \6624 , \6625 ,         \6626 , \6627 , \6628 , \6629 , \6630 , \6631 , \6632 , \6633 , \6634 , \6635 ,         \6636 , \6637 , \6638 , \6639 , \6640 , \6641 , \6642 , \6643 , \6644 , \6645 ,         \6646 , \6647 , \6648 , \6649 , \6650 , \6651 , \6652 , \6653 , \6654 , \6655 ,         \6656 , \6657 , \6658 , \6659 , \6660 , \6661 , \6662 , \6663 , \6664 , \6665 ,         \6666 , \6667 , \6668 , \6669 , \6670 , \6671 , \6672 , \6673 , \6674 , \6675 ,         \6676 , \6677 , \6678 , \6679 , \6680 , \6681 , \6682 , \6683 , \6684 , \6685 ,         \6686 , \6687 , \6688 , \6689 , \6690 , \6691 , \6692 , \6693 , \6694 , \6695 ,         \6696 , \6697 , \6698 , \6699 , \6700 , \6701 , \6702 , \6703 , \6704 , \6705 ,         \6706 , \6707 , \6708 , \6709 , \6710 , \6711 , \6712 , \6713 , \6714 , \6715 ,         \6716 , \6717 , \6718 , \6719 , \6720 , \6721 , \6722 , \6723 , \6724 , \6725 ,         \6726 , \6727 , \6728 , \6729 , \6730 , \6731 , \6732 , \6733 , \6734 , \6735 ,         \6736 , \6737 , \6738 , \6739 , \6740 , \6741 , \6742 , \6743 , \6744 , \6745 ,         \6746 , \6747 , \6748 , \6749 , \6750 , \6751 , \6752 , \6753 , \6754 , \6755 ,         \6756 , \6757 , \6758 , \6759 , \6760 , \6761 , \6762 , \6763 , \6764 , \6765 ,         \6766 , \6767 , \6768 , \6769 , \6770 , \6771 , \6772 , \6773 , \6774 , \6775 ,         \6776 , \6777 , \6778 , \6779 , \6780 , \6781 , \6782 , \6783 , \6784 , \6785 ,         \6786 , \6787 , \6788 , \6789 , \6790 , \6791 , \6792 , \6793 , \6794 , \6795 ,         \6796 , \6797 , \6798 , \6799 , \6800 , \6801 , \6802 , \6803 , \6804 , \6805 ,         \6806 , \6807 , \6808 , \6809 , \6810 , \6811 , \6812 , \6813 , \6814 , \6815 ,         \6816 , \6817 , \6818 , \6819 , \6820 , \6821 , \6822 , \6823 , \6824 , \6825 ,         \6826 , \6827 , \6828 , \6829 , \6830 , \6831 , \6832 , \6833 , \6834 , \6835 ,         \6836 , \6837 , \6838 , \6839 , \6840 , \6841 , \6842 , \6843 , \6844 , \6845 ,         \6846 , \6847 , \6848 , \6849 , \6850 , \6851 , \6852 , \6853 , \6854 , \6855 ,         \6856 , \6857 , \6858 , \6859 , \6860 , \6861 , \6862 , \6863 , \6864 , \6865 ,         \6866 , \6867 , \6868 , \6869 , \6870 , \6871 , \6872 , \6873 , \6874 , \6875 ,         \6876 , \6877 , \6878 , \6879 , \6880 , \6881 , \6882 , \6883 , \6884 , \6885 ,         \6886 , \6887 , \6888 , \6889 , \6890 , \6891 , \6892 , \6893 , \6894 , \6895 ,         \6896 , \6897 , \6898 , \6899 , \6900 , \6901 , \6902 , \6903 , \6904 , \6905 ,         \6906 , \6907 , \6908 , \6909 , \6910 , \6911 , \6912 , \6913 , \6914 , \6915 ,         \6916 , \6917 , \6918 , \6919 , \6920 , \6921 , \6922 , \6923 , \6924 , \6925 ,         \6926 , \6927 , \6928 , \6929 , \6930 , \6931 , \6932 , \6933 , \6934 , \6935 ,         \6936 , \6937 , \6938 , \6939 , \6940 , \6941 , \6942 , \6943 , \6944 , \6945 ,         \6946 , \6947 , \6948 , \6949 , \6950 , \6951 , \6952 , \6953 , \6954 , \6955 ,         \6956 , \6957 , \6958 , \6959 , \6960 , \6961 , \6962 , \6963 , \6964 , \6965 ,         \6966 , \6967 , \6968 , \6969 , \6970 , \6971 , \6972 , \6973 , \6974 , \6975 ,         \6976 , \6977 , \6978 , \6979 , \6980 , \6981 , \6982 , \6983 , \6984 , \6985 ,         \6986 , \6987 , \6988 , \6989 , \6990 , \6991 , \6992 , \6993 , \6994 , \6995 ,         \6996 , \6997 , \6998 , \6999 , \7000 , \7001 , \7002 , \7003 , \7004 , \7005 ,         \7006 , \7007 , \7008 , \7009 , \7010 , \7011 , \7012 , \7013 , \7014 , \7015 ,         \7016 , \7017 , \7018 , \7019 , \7020 , \7021 , \7022 , \7023 , \7024 , \7025 ,         \7026 , \7027 , \7028 , \7029 , \7030 , \7031 , \7032 , \7033 , \7034 , \7035 ,         \7036 , \7037 , \7038 , \7039 , \7040 , \7041 , \7042 , \7043 , \7044 , \7045 ,         \7046 , \7047 , \7048 , \7049 , \7050 , \7051 , \7052 , \7053 , \7054 , \7055 ,         \7056 , \7057 , \7058 , \7059 , \7060 , \7061 , \7062 , \7063 , \7064 , \7065 ,         \7066 , \7067 , \7068 , \7069 , \7070 , \7071 , \7072 , \7073 , \7074 , \7075 ,         \7076 , \7077 , \7078 , \7079 , \7080 , \7081 , \7082 , \7083 , \7084 , \7085 ,         \7086 , \7087 , \7088 , \7089 , \7090 , \7091 , \7092 , \7093 , \7094 , \7095 ,         \7096 , \7097 , \7098 , \7099 , \7100 , \7101 , \7102 , \7103 , \7104 , \7105 ,         \7106 , \7107 , \7108 , \7109 , \7110 , \7111 , \7112 , \7113 , \7114 , \7115 ,         \7116 , \7117 , \7118 , \7119 , \7120 , \7121 , \7122 , \7123 , \7124 , \7125 ,         \7126 , \7127 , \7128 , \7129 , \7130 , \7131 , \7132 , \7133 , \7134 , \7135 ,         \7136 , \7137 , \7138 , \7139 , \7140 , \7141 , \7142 , \7143 , \7144 , \7145 ,         \7146 , \7147 , \7148 , \7149 , \7150 , \7151 , \7152 , \7153 , \7154 , \7155 ,         \7156 , \7157 , \7158 , \7159 , \7160 , \7161 , \7162 , \7163 , \7164 , \7165 ,         \7166 , \7167 , \7168 , \7169 , \7170 , \7171 , \7172 , \7173 , \7174 , \7175 ,         \7176 , \7177 , \7178 , \7179 , \7180 , \7181 , \7182 , \7183 , \7184 , \7185 ,         \7186 , \7187 , \7188 , \7189 , \7190 , \7191 , \7192 , \7193 , \7194 , \7195 ,         \7196 , \7197 , \7198 , \7199 , \7200 , \7201 , \7202 , \7203 , \7204 , \7205 ,         \7206 , \7207 , \7208 , \7209 , \7210 , \7211 , \7212 , \7213 , \7214 , \7215 ,         \7216 , \7217 , \7218 , \7219 , \7220 , \7221 , \7222 , \7223 , \7224 , \7225 ,         \7226 , \7227 , \7228 , \7229 , \7230 , \7231 , \7232 , \7233 , \7234 , \7235 ,         \7236 , \7237 , \7238 , \7239 , \7240 , \7241 , \7242 , \7243 , \7244 , \7245 ,         \7246 , \7247 , \7248 , \7249 , \7250 , \7251 , \7252 , \7253 , \7254 , \7255 ,         \7256 , \7257 , \7258 , \7259 , \7260 , \7261 , \7262 , \7263 , \7264 , \7265 ,         \7266 , \7267 , \7268 , \7269 , \7270 , \7271 , \7272 , \7273 , \7274 , \7275 ,         \7276 , \7277 , \7278 , \7279 , \7280 , \7281 , \7282 , \7283 , \7284 , \7285 ,         \7286 , \7287 , \7288 , \7289 , \7290 , \7291 , \7292 , \7293 , \7294 , \7295 ,         \7296 , \7297 , \7298 , \7299 , \7300 , \7301 , \7302 , \7303 , \7304 , \7305 ,         \7306 , \7307 , \7308 , \7309 , \7310 , \7311 , \7312 , \7313 , \7314 , \7315 ,         \7316 , \7317 , \7318 , \7319 , \7320 , \7321 , \7322 , \7323 , \7324 , \7325 ,         \7326 , \7327 , \7328 , \7329 , \7330 , \7331 , \7332 , \7333 , \7334 , \7335 ,         \7336 , \7337 , \7338 , \7339 , \7340 , \7341 , \7342 , \7343 , \7344 , \7345 ,         \7346 , \7347 , \7348 , \7349 , \7350 , \7351 , \7352 , \7353 , \7354 , \7355 ,         \7356 , \7357 , \7358 , \7359 , \7360 , \7361 , \7362 , \7363 , \7364 , \7365 ,         \7366 , \7367 , \7368 , \7369 , \7370 , \7371 , \7372 , \7373 , \7374 , \7375 ,         \7376 , \7377 , \7378 , \7379 , \7380 , \7381 , \7382 , \7383 , \7384 , \7385 ,         \7386 , \7387 , \7388 , \7389 , \7390 , \7391 , \7392 , \7393 , \7394 , \7395 ,         \7396 , \7397 , \7398 , \7399 , \7400 , \7401 , \7402 , \7403 , \7404 , \7405 ,         \7406 , \7407 , \7408 , \7409 , \7410 , \7411 , \7412 , \7413 , \7414 , \7415 ,         \7416 , \7417 , \7418 , \7419 , \7420 , \7421 , \7422 , \7423 , \7424 , \7425 ,         \7426 , \7427 , \7428 , \7429 , \7430 , \7431 , \7432 , \7433 , \7434 , \7435 ,         \7436 , \7437 , \7438 , \7439 , \7440 , \7441 , \7442 , \7443 , \7444 , \7445 ,         \7446 , \7447 , \7448 , \7449 , \7450 , \7451 , \7452 , \7453 , \7454 , \7455 ,         \7456 , \7457 , \7458 , \7459 , \7460 , \7461 , \7462 , \7463 , \7464 , \7465 ,         \7466 , \7467 , \7468 , \7469 , \7470 , \7471 , \7472 , \7473 , \7474 , \7475 ,         \7476 , \7477 , \7478 , \7479 , \7480 , \7481 , \7482 , \7483 , \7484 , \7485 ,         \7486 , \7487 , \7488 , \7489 , \7490 , \7491 , \7492 , \7493 , \7494 , \7495 ,         \7496 , \7497 , \7498 , \7499 , \7500 , \7501 , \7502 , \7503 , \7504 , \7505 ,         \7506 , \7507 , \7508 ;
mbuf \U$labaj768 ( \o[31] , \7238 );
mbuf \U$labaj769 ( \o[30] , \7251 );
mbuf \U$labaj770 ( \o[29] , \7262 );
mbuf \U$labaj771 ( \o[28] , \7274 );
mbuf \U$labaj772 ( \o[27] , \7288 );
mbuf \U$labaj773 ( \o[26] , \7300 );
mbuf \U$labaj774 ( \o[25] , \7311 );
mbuf \U$labaj775 ( \o[24] , \7343 );
mbuf \U$labaj776 ( \o[23] , \7337 );
mbuf \U$labaj777 ( \o[22] , \7508 );
mbuf \U$labaj778 ( \o[21] , \7354 );
mbuf \U$labaj779 ( \o[20] , \7360 );
mbuf \U$labaj780 ( \o[19] , \7375 );
mbuf \U$labaj781 ( \o[18] , \7381 );
mbuf \U$labaj782 ( \o[17] , \7392 );
mbuf \U$labaj783 ( \o[16] , \7398 );
mbuf \U$labaj784 ( \o[15] , \7418 );
mbuf \U$labaj785 ( \o[14] , \7426 );
mbuf \U$labaj786 ( \o[13] , \7436 );
mbuf \U$labaj787 ( \o[12] , \7458 );
mbuf \U$labaj788 ( \o[11] , \7452 );
mbuf \U$labaj789 ( \o[10] , \7464 );
mbuf \U$labaj790 ( \o[9] , \7474 );
mbuf \U$labaj791 ( \o[8] , \7480 );
mbuf \U$labaj792 ( \o[7] , \7482 );
mbuf \U$labaj793 ( \o[6] , \7507 );
mbuf \U$labaj794 ( \o[5] , \7488 );
mbuf \U$labaj795 ( \o[4] , \7495 );
mbuf \U$labaj796 ( \o[3] , \7497 );
mbuf \U$labaj797 ( \o[2] , \7502 );
mbuf \U$labaj798 ( \o[1] , \7505 );
mbuf \U$labaj799 ( \o[0] , \7506 );
mnot \g4514/U$3 ( \99 , \d[15] );
mxor \g36663/U$1 ( \100 , \b[3] , \a[2] );
mnot \mul_6_11_g6696/U$3 ( \101 , \100 );
mxnor \mul_6_11_g6910/U$1 ( \102 , \b[3] , \b[2] );
mxor \mul_6_11_g36689/U$1 ( \103 , \b[2] , \b[1] );
mnor \mul_6_11_g6763/U$1 ( \104 , \102 , \103 );
mnot \mul_6_11_g6696/U$4 ( \105 , \104 );
mor \mul_6_11_g6696/U$2 ( \106 , \101 , \105 );
mxor \g36662/U$1 ( \107 , \b[3] , \a[3] );
mnand \mul_6_11_g6747/U$1 ( \108 , \103 , \107 );
mnand \mul_6_11_g6696/U$1 ( \109 , \106 , \108 );
mor \mul_6_11_g6803/U$2 ( \110 , \a[0] , \b[4] );
mnand \mul_6_11_g6803/U$1 ( \111 , \110 , \b[3] );
mnand \mul_6_11_g6880/U$1 ( \112 , \a[0] , \b[4] );
mnand \mul_6_11_g6786/U$1 ( \113 , \111 , \112 , \b[5] );
mnot \mul_6_11_g6785/U$1 ( \114 , \113 );
mand \mul_6_11_g6661/U$1 ( \115 , \109 , \114 );
mnot \mul_6_11_g6922/U$2 ( \116 , \115 );
mxor \mul_6_11_g6840/U$1 ( \117 , \a[5] , \b[1] );
mnot \mul_6_11_g6733/U$3 ( \118 , \117 );
mnot \mul_6_11_g6899/U$2 ( \119 , \b[1] );
mnor \mul_6_11_g6899/U$1 ( \120 , \119 , \b[0] );
mnot \mul_6_11_g6733/U$4 ( \121 , \120 );
mor \mul_6_11_g6733/U$2 ( \122 , \118 , \121 );
mxor \mul_6_11_g6817/U$1 ( \123 , \a[6] , \b[1] );
mnand \mul_6_11_g6750/U$1 ( \124 , \123 , \b[0] );
mnand \mul_6_11_g6733/U$1 ( \125 , \122 , \124 );
mnot \mul_6_11_g6732/U$1 ( \126 , \125 );
mnand \mul_6_11_g6922/U$1 ( \127 , \116 , \126 );
mnot \mul_6_11_g6580/U$3 ( \128 , \127 );
mxor \mul_6_11_g36836/U$1 ( \129 , \b[6] , \b[5] );
mand \g37047/U$1 ( \130 , \129 , \a[0] );
mxor \mul_6_11_g6862/U$1 ( \131 , \a[1] , \b[5] );
mnot \mul_6_11_g6665/U$3 ( \132 , \131 );
mxor \mul_6_11_g6903/U$1 ( \133 , \b[5] , \b[4] );
mnot \mul_6_11_g6714/U$2 ( \134 , \133 );
mxor \mul_6_11_g36679/U$1 ( \135 , \b[4] , \b[3] );
mnor \mul_6_11_g6714/U$1 ( \136 , \134 , \135 );
mnot \mul_6_11_g6665/U$4 ( \137 , \136 );
mor \mul_6_11_g6665/U$2 ( \138 , \132 , \137 );
mxor \mul_6_11_g36677/U$1 ( \139 , \b[4] , \b[3] );
mxor \mul_6_11_g6855/U$1 ( \140 , \a[2] , \b[5] );
mnand \mul_6_11_g6709/U$1 ( \141 , \139 , \140 );
mnand \mul_6_11_g6665/U$1 ( \142 , \138 , \141 );
mxor \mul_6_11_g6613/U$1 ( \143 , \130 , \142 );
mnot \mul_6_11_g6698/U$3 ( \144 , \107 );
mnot \mul_6_11_g6698/U$4 ( \145 , \104 );
mor \mul_6_11_g6698/U$2 ( \146 , \144 , \145 );
mxor \mul_6_11_g36681/U$1 ( \147 , \b[2] , \b[1] );
mxor \mul_6_11_g6837/U$1 ( \148 , \a[4] , \b[3] );
mnand \mul_6_11_g6753/U$1 ( \149 , \147 , \148 );
mnand \mul_6_11_g6698/U$1 ( \150 , \146 , \149 );
mxor \mul_6_11_g6613/U$1_r1 ( \151 , \143 , \150 );
mnot \mul_6_11_g6580/U$4 ( \152 , \151 );
mor \mul_6_11_g6580/U$2 ( \153 , \128 , \152 );
mnand \mul_6_11_g6629/U$1 ( \154 , \115 , \125 );
mnand \mul_6_11_g6580/U$1 ( \155 , \153 , \154 );
mor \mul_6_11_g6801/U$2 ( \156 , \a[0] , \b[6] );
mnand \mul_6_11_g6801/U$1 ( \157 , \156 , \b[5] );
mnand \mul_6_11_g6874/U$1 ( \158 , \a[0] , \b[6] );
mnand \mul_6_11_g6789/U$1 ( \159 , \157 , \158 , \b[7] );
mnot \mul_6_11_g6652/U$3 ( \160 , \159 );
mnot \mul_6_11_g6699/U$3 ( \161 , \148 );
mnot \mul_6_11_g6699/U$4 ( \162 , \104 );
mor \mul_6_11_g6699/U$2 ( \163 , \161 , \162 );
mxor \g36661/U$1 ( \164 , \b[3] , \a[5] );
mnand \mul_6_11_g6755/U$1 ( \165 , \147 , \164 );
mnand \mul_6_11_g6699/U$1 ( \166 , \163 , \165 );
mnot \mul_6_11_g6652/U$4 ( \167 , \166 );
mor \mul_6_11_g6652/U$2 ( \168 , \160 , \167 );
mor \mul_6_11_g6652/U$5 ( \169 , \166 , \159 );
mnand \mul_6_11_g6652/U$1 ( \170 , \168 , \169 );
mxor \mul_6_11_g6613/U$4 ( \171 , \130 , \142 );
mand \mul_6_11_g6613/U$3 ( \172 , \171 , \150 );
mand \mul_6_11_g6613/U$5 ( \173 , \130 , \142 );
mor \mul_6_11_g6613/U$2 ( \174 , \172 , \173 );
mxor \mul_6_11_g6549/U$1 ( \175 , \170 , \174 );
mnot \mul_6_11_g6734/U$3 ( \176 , \123 );
mnot \mul_6_11_g6734/U$4 ( \177 , \120 );
mor \mul_6_11_g6734/U$2 ( \178 , \176 , \177 );
mxor \mul_6_11_g6824/U$1 ( \179 , \a[7] , \b[1] );
mnand \mul_6_11_g6756/U$1 ( \180 , \179 , \b[0] );
mnand \mul_6_11_g6734/U$1 ( \181 , \178 , \180 );
mxor \mul_6_11_g6867/U$1 ( \182 , \a[0] , \b[7] );
mnot \mul_6_11_g6690/U$3 ( \183 , \182 );
mxor \mul_6_11_g6829/U$1 ( \184 , \b[6] , \b[5] );
mxnor \mul_6_11_g6909/U$1 ( \185 , \b[7] , \b[6] );
mnor \mul_6_11_g6794/U$1 ( \186 , \184 , \185 );
mnot \mul_6_11_g6690/U$4 ( \187 , \186 );
mor \mul_6_11_g6690/U$2 ( \188 , \183 , \187 );
mxor \g36666/U$1 ( \189 , \b[7] , \a[1] );
mnand \mul_6_11_g6757/U$1 ( \190 , \129 , \189 );
mnand \mul_6_11_g6690/U$1 ( \191 , \188 , \190 );
mxor \mul_6_11_g6618/U$1 ( \192 , \181 , \191 );
mnot \mul_6_11_g6666/U$3 ( \193 , \140 );
mnot \mul_6_11_g6715/U$2 ( \194 , \133 );
mnor \mul_6_11_g6715/U$1 ( \195 , \194 , \135 );
mnot \mul_6_11_g6666/U$4 ( \196 , \195 );
mor \mul_6_11_g6666/U$2 ( \197 , \193 , \196 );
mxor \mul_6_11_g6854/U$1 ( \198 , \a[3] , \b[5] );
mnand \mul_6_11_g6710/U$1 ( \199 , \139 , \198 );
mnand \mul_6_11_g6666/U$1 ( \200 , \197 , \199 );
mxor \mul_6_11_g6618/U$1_r1 ( \201 , \192 , \200 );
mxor \mul_6_11_g6549/U$1_r1 ( \202 , \175 , \201 );
mxor \mul_6_11_g6500/U$4 ( \203 , \155 , \202 );
mnot \mul_6_11_g6695/U$1 ( \204 , \109 );
mxnor \g36659/U$1 ( \205 , \204 , \113 );
mnot \mul_6_11_g6839/U$1 ( \206 , \117 );
mnot \g37080/U$3 ( \207 , \206 );
mnot \mul_6_11_g6902/U$1 ( \208 , \b[0] );
mnot \g37080/U$4 ( \209 , \208 );
mand \g37080/U$2 ( \210 , \207 , \209 );
mnot \mul_6_11_g6898/U$2 ( \211 , \b[1] );
mnor \mul_6_11_g6898/U$1 ( \212 , \211 , \b[0] );
mxor \mul_6_11_g6841/U$1 ( \213 , \a[4] , \b[1] );
mand \g37080/U$5 ( \214 , \212 , \213 );
mnor \g37080/U$1 ( \215 , \210 , \214 );
mxor \mul_6_11_g36755/U$1 ( \216 , \a[0] , \b[5] );
mnor \mul_6_11_g6881/U$1 ( \217 , \b[4] , \b[3] );
mnand \mul_6_11_g6680/U$1 ( \218 , \216 , \133 , \217 );
mand \mul_6_11_g6907/U$1 ( \219 , \b[4] , \b[3] );
mnand \mul_6_11_g6679/U$1 ( \220 , \216 , \133 , \219 );
mnand \mul_6_11_g6711/U$1 ( \221 , \135 , \131 );
mand \mul_6_11_g6654/U$1 ( \222 , \218 , \220 , \221 );
mand \mul_6_11_g6614/U$2 ( \223 , \215 , \222 );
mor \mul_6_11_g6587/U$2 ( \224 , \205 , \223 );
mor \mul_6_11_g6924/U$1 ( \225 , \222 , \215 );
mnand \mul_6_11_g6587/U$1 ( \226 , \224 , \225 );
mnot \mul_6_11_g6558/U$2 ( \227 , \226 );
mnot \mul_6_11_g6581/U$3 ( \228 , \151 );
mand \mul_6_11_g6660/U$1 ( \229 , \109 , \114 );
mnot \mul_6_11_g6609/U$3 ( \230 , \229 );
mnot \mul_6_11_g6609/U$4 ( \231 , \126 );
mand \mul_6_11_g6609/U$2 ( \232 , \230 , \231 );
mand \mul_6_11_g6609/U$5 ( \233 , \115 , \126 );
mnor \mul_6_11_g6609/U$1 ( \234 , \232 , \233 );
mnot \mul_6_11_g6581/U$4 ( \235 , \234 );
mand \mul_6_11_g6581/U$2 ( \236 , \228 , \235 );
mand \mul_6_11_g6581/U$5 ( \237 , \151 , \234 );
mnor \mul_6_11_g6581/U$1 ( \238 , \236 , \237 );
mnand \mul_6_11_g6558/U$1 ( \239 , \227 , \238 );
mnot \g36749/U$3 ( \240 , \239 );
mnand \mul_6_11_g6718/U$1 ( \241 , \139 , \a[0] );
mnot \mul_6_11_g6643/U$3 ( \242 , \241 );
mxor \mul_6_11_g6852/U$1 ( \243 , \a[3] , \b[1] );
mnot \mul_6_11_g6739/U$3 ( \244 , \243 );
mnot \mul_6_11_g6739/U$4 ( \245 , \212 );
mor \mul_6_11_g6739/U$2 ( \246 , \244 , \245 );
mnand \mul_6_11_g6769/U$1 ( \247 , \213 , \b[0] );
mnand \mul_6_11_g6739/U$1 ( \248 , \246 , \247 );
mnot \mul_6_11_g6738/U$1 ( \249 , \248 );
mnot \mul_6_11_g6643/U$4 ( \250 , \249 );
mor \mul_6_11_g6643/U$2 ( \251 , \242 , \250 );
mxor \mul_6_11_g6856/U$1 ( \252 , \a[1] , \b[3] );
mnot \mul_6_11_g6702/U$3 ( \253 , \252 );
mnot \mul_6_11_g6702/U$4 ( \254 , \104 );
mor \mul_6_11_g6702/U$2 ( \255 , \253 , \254 );
mnand \mul_6_11_g6754/U$1 ( \256 , \147 , \100 );
mnand \mul_6_11_g6702/U$1 ( \257 , \255 , \256 );
mnand \mul_6_11_g6643/U$1 ( \258 , \251 , \257 );
mnot \mul_6_11_g6926/U$2 ( \259 , \241 );
mnand \mul_6_11_g6926/U$1 ( \260 , \259 , \248 );
mnand \mul_6_11_g6631/U$1 ( \261 , \258 , \260 );
mnot \mul_6_11_g6622/U$1 ( \262 , \261 );
mnot \mul_6_11_g6545/U$3 ( \263 , \262 );
mxor \mul_6_11_g6593/U$1 ( \264 , \113 , \204 );
mxor \mul_6_11_g6614/U$1 ( \265 , \215 , \222 );
mxnor \mul_6_11_g6593/U$1_r1 ( \266 , \264 , \265 );
mnot \mul_6_11_g6545/U$4 ( \267 , \266 );
mor \mul_6_11_g6545/U$2 ( \268 , \263 , \267 );
mand \g36745/U$2 ( \269 , \248 , \241 );
mnot \g36745/U$4 ( \270 , \248 );
mand \g36746/U$1 ( \271 , \139 , \a[0] );
mand \g36745/U$3 ( \272 , \270 , \271 );
mnor \g36745/U$1 ( \273 , \269 , \272 );
mand \mul_6_11_g6633/U$2 ( \274 , \273 , \257 );
mnot \mul_6_11_g6633/U$4 ( \275 , \273 );
mnot \mul_6_11_g6701/U$1 ( \276 , \257 );
mand \mul_6_11_g6633/U$3 ( \277 , \275 , \276 );
mnor \mul_6_11_g6633/U$1 ( \278 , \274 , \277 );
mnand \mul_6_11_g6879/U$1 ( \279 , \a[0] , \b[2] );
mor \mul_6_11_g6802/U$2 ( \280 , \a[0] , \b[2] );
mnand \mul_6_11_g6802/U$1 ( \281 , \280 , \b[1] );
mnand \g37136/U$1 ( \282 , \279 , \b[3] , \281 );
mnot \mul_6_11_g6928/U$2 ( \283 , \282 );
mxor \mul_6_11_g6851/U$1 ( \284 , \a[2] , \b[1] );
mnot \mul_6_11_g6741/U$3 ( \285 , \284 );
mnot \mul_6_11_g6741/U$4 ( \286 , \212 );
mor \mul_6_11_g6741/U$2 ( \287 , \285 , \286 );
mnand \mul_6_11_g6767/U$1 ( \288 , \243 , \b[0] );
mnand \mul_6_11_g6741/U$1 ( \289 , \287 , \288 );
mnand \mul_6_11_g6928/U$1 ( \290 , \283 , \289 );
mnand \mul_6_11_g6597/U$1 ( \291 , \278 , \290 );
mnot \g37134/U$3 ( \292 , \291 );
mxor \g36667/U$1 ( \293 , \b[3] , \a[0] );
mnot \mul_6_11_g6704/U$3 ( \294 , \293 );
mnor \mul_6_11_g6764/U$1 ( \295 , \102 , \103 );
mnot \mul_6_11_g6704/U$4 ( \296 , \295 );
mor \mul_6_11_g6704/U$2 ( \297 , \294 , \296 );
mnand \mul_6_11_g6751/U$1 ( \298 , \147 , \252 );
mnand \mul_6_11_g6704/U$1 ( \299 , \297 , \298 );
mnot \mul_6_11_g6641/U$2 ( \300 , \299 );
mxor \g36673/U$1 ( \301 , \289 , \282 );
mnand \mul_6_11_g6641/U$1 ( \302 , \300 , \301 );
mnot \g37135/U$3 ( \303 , \302 );
mnand \mul_6_11_g6779/U$1 ( \304 , \147 , \a[0] );
mnot \g37079/U$2 ( \305 , \304 );
mxor \g36664/U$1 ( \306 , \b[1] , \a[1] );
mnot \mul_6_11_g6742/U$3 ( \307 , \306 );
mnot \mul_6_11_g6742/U$4 ( \308 , \120 );
mor \mul_6_11_g6742/U$2 ( \309 , \307 , \308 );
mnand \mul_6_11_g6768/U$1 ( \310 , \284 , \b[0] );
mnand \mul_6_11_g6742/U$1 ( \311 , \309 , \310 );
mnor \g37079/U$1 ( \312 , \305 , \311 );
mnot \mul_6_11_g6723/U$3 ( \313 , \b[0] );
mnot \mul_6_11_g6857/U$1 ( \314 , \306 );
mnot \mul_6_11_g6723/U$4 ( \315 , \314 );
mor \mul_6_11_g6723/U$2 ( \316 , \313 , \315 );
mnand \mul_6_11_g6883/U$1 ( \317 , \a[0] , \b[0] );
mnand \mul_6_11_g6806/U$1 ( \318 , \317 , \b[1] );
mnor \mul_6_11_g6773/U$1 ( \319 , \318 , \a[0] );
mnand \mul_6_11_g6723/U$1 ( \320 , \316 , \319 );
mor \mul_6_11_g6648/U$2 ( \321 , \312 , \320 );
mnot \g36921/U$2 ( \322 , \304 );
mnand \g36921/U$1 ( \323 , \322 , \311 );
mnand \mul_6_11_g6648/U$1 ( \324 , \321 , \323 );
mnot \g37135/U$4 ( \325 , \324 );
mor \g37135/U$2 ( \326 , \303 , \325 );
mnot \mul_6_11_g6925/U$2 ( \327 , \301 );
mnand \mul_6_11_g6925/U$1 ( \328 , \327 , \299 );
mnand \g37135/U$1 ( \329 , \326 , \328 );
mnot \g37134/U$4 ( \330 , \329 );
mor \g37134/U$2 ( \331 , \292 , \330 );
mnot \mul_6_11_g6619/U$1 ( \332 , \278 );
mnot \mul_6_11_g6657/U$1 ( \333 , \290 );
mnand \mul_6_11_g6595/U$1 ( \334 , \332 , \333 );
mnand \g37134/U$1 ( \335 , \331 , \334 );
mnand \mul_6_11_g6545/U$1 ( \336 , \268 , \335 );
mnot \fopt36949/U$1 ( \337 , \266 );
mnand \mul_6_11_g6570/U$1 ( \338 , \337 , \261 );
mnand \mul_6_11_g6539/U$1 ( \339 , \336 , \338 );
mnot \g36749/U$4 ( \340 , \339 );
mor \g36749/U$2 ( \341 , \240 , \340 );
mnot \mul_6_11_g6919/U$2 ( \342 , \238 );
mnand \mul_6_11_g6919/U$1 ( \343 , \342 , \226 );
mnand \g36749/U$1 ( \344 , \341 , \343 );
mand \mul_6_11_g6500/U$3 ( \345 , \203 , \344 );
mand \mul_6_11_g6500/U$5 ( \346 , \155 , \202 );
mor \mul_6_11_g6500/U$2 ( \347 , \345 , \346 );
mnot \mul_6_11_g6726/U$3 ( \348 , \120 );
mxor \mul_6_11_g36904/U$1 ( \349 , \a[8] , \b[1] );
mnot \mul_6_11_g6726/U$4 ( \350 , \349 );
mor \mul_6_11_g6726/U$2 ( \351 , \348 , \350 );
mxor \mul_6_11_g6825/U$1 ( \352 , \a[9] , \b[1] );
mnand \mul_6_11_g6772/U$1 ( \353 , \352 , \b[0] );
mnand \mul_6_11_g6726/U$1 ( \354 , \351 , \353 );
mxor \g36665/U$1 ( \355 , \b[7] , \a[2] );
mnot \mul_6_11_g6689/U$3 ( \356 , \355 );
mnot \mul_6_11_g6689/U$4 ( \357 , \186 );
mor \mul_6_11_g6689/U$2 ( \358 , \356 , \357 );
mxor \mul_6_11_g37179/U$1 ( \359 , \a[3] , \b[7] );
mnand \mul_6_11_g37183/U$1 ( \360 , \359 , \129 );
mnand \mul_6_11_g6689/U$1 ( \361 , \358 , \360 );
mxor \mul_6_11_g6627/U$1 ( \362 , \354 , \361 );
mxor \mul_6_11_g6811/U$1 ( \363 , \a[6] , \b[3] );
mnot \mul_6_11_g6697/U$3 ( \364 , \363 );
mnot \mul_6_11_g6697/U$4 ( \365 , \295 );
mor \mul_6_11_g6697/U$2 ( \366 , \364 , \365 );
mxor \mul_6_11_g6812/U$1 ( \367 , \a[7] , \b[3] );
mnand \mul_6_11_g6746/U$1 ( \368 , \147 , \367 );
mnand \mul_6_11_g6697/U$1 ( \369 , \366 , \368 );
mxor \mul_6_11_g6627/U$1_r1 ( \370 , \362 , \369 );
mnot \fopt36722/U$1 ( \371 , \370 );
mnot \mul_6_11_g6577/U$3 ( \372 , \371 );
mnot \mul_6_11_g6688/U$3 ( \373 , \189 );
mnor \mul_6_11_g6795/U$1 ( \374 , \185 , \184 );
mnot \mul_6_11_g6688/U$4 ( \375 , \374 );
mor \mul_6_11_g6688/U$2 ( \376 , \373 , \375 );
mnand \mul_6_11_g6748/U$1 ( \377 , \129 , \355 );
mnand \mul_6_11_g6688/U$1 ( \378 , \376 , \377 );
mnot \mul_6_11_g6663/U$3 ( \379 , \198 );
mnot \mul_6_11_g6663/U$4 ( \380 , \195 );
mor \mul_6_11_g6663/U$2 ( \381 , \379 , \380 );
mxor \mul_6_11_g37180/U$1 ( \382 , \a[4] , \b[5] );
mnand \mul_6_11_g6708/U$1 ( \383 , \139 , \382 );
mnand \mul_6_11_g6663/U$1 ( \384 , \381 , \383 );
mxor \mul_6_11_g6591/U$4 ( \385 , \378 , \384 );
mnot \mul_6_11_g2/U$2 ( \386 , \166 );
mnor \mul_6_11_g2/U$1 ( \387 , \386 , \159 );
mand \mul_6_11_g6591/U$3 ( \388 , \385 , \387 );
mand \mul_6_11_g6591/U$5 ( \389 , \378 , \384 );
mor \mul_6_11_g6591/U$2 ( \390 , \388 , \389 );
mnot \mul_6_11_g6577/U$4 ( \391 , \390 );
mor \mul_6_11_g6577/U$2 ( \392 , \372 , \391 );
mnot \fopt36723/U$1 ( \393 , \370 );
mor \mul_6_11_g6577/U$5 ( \394 , \393 , \390 );
mnand \mul_6_11_g6577/U$1 ( \395 , \392 , \394 );
mnot \mul_6_11_g6542/U$3 ( \396 , \395 );
mxor \mul_6_11_g6863/U$1 ( \397 , \a[0] , \b[9] );
mnot \mul_6_11_g6684/U$3 ( \398 , \397 );
mxnor \g37137/U$1 ( \399 , \b[9] , \b[8] );
mxor \mul_6_11_g36686/U$1 ( \400 , \b[8] , \b[7] );
mnor \mul_6_11_g6796/U$1 ( \401 , \399 , \400 );
mnot \mul_6_11_g6684/U$4 ( \402 , \401 );
mor \mul_6_11_g6684/U$2 ( \403 , \398 , \402 );
mxor \mul_6_11_g6868/U$1 ( \404 , \a[1] , \b[9] );
mnand \mul_6_11_g6752/U$1 ( \405 , \400 , \404 );
mnand \mul_6_11_g6684/U$1 ( \406 , \403 , \405 );
mnot \fopt36882/U$1 ( \407 , \406 );
mnot \mul_6_11_g6601/U$3 ( \408 , \407 );
mor \mul_6_11_g6800/U$2 ( \409 , \a[0] , \b[8] );
mnand \mul_6_11_g6800/U$1 ( \410 , \409 , \b[7] );
mnand \mul_6_11_g6871/U$1 ( \411 , \a[0] , \b[8] );
mand \mul_6_11_g6906/U$1 ( \412 , \410 , \411 , \b[9] );
mnot \mul_6_11_g6664/U$3 ( \413 , \382 );
mnot \mul_6_11_g6664/U$4 ( \414 , \136 );
mor \mul_6_11_g6664/U$2 ( \415 , \413 , \414 );
mxor \mul_6_11_g37181/U$1 ( \416 , \a[5] , \b[5] );
mnand \mul_6_11_g6707/U$1 ( \417 , \139 , \416 );
mnand \mul_6_11_g6664/U$1 ( \418 , \415 , \417 );
mxor \mul_6_11_g6635/U$1 ( \419 , \412 , \418 );
mnot \mul_6_11_g6601/U$4 ( \420 , \419 );
mor \mul_6_11_g6601/U$2 ( \421 , \408 , \420 );
mor \mul_6_11_g6601/U$5 ( \422 , \419 , \407 );
mnand \mul_6_11_g6601/U$1 ( \423 , \421 , \422 );
mand \mul_6_11_g6770/U$1 ( \424 , \400 , \a[0] );
mnot \mul_6_11_g6728/U$3 ( \425 , \179 );
mnot \mul_6_11_g6728/U$4 ( \426 , \120 );
mor \mul_6_11_g6728/U$2 ( \427 , \425 , \426 );
mnand \mul_6_11_g6775/U$1 ( \428 , \349 , \b[0] );
mnand \mul_6_11_g6728/U$1 ( \429 , \427 , \428 );
mxor \mul_6_11_g6612/U$4 ( \430 , \424 , \429 );
mnot \mul_6_11_g6700/U$3 ( \431 , \164 );
mnot \mul_6_11_g6700/U$4 ( \432 , \295 );
mor \mul_6_11_g6700/U$2 ( \433 , \431 , \432 );
mnand \mul_6_11_g6758/U$1 ( \434 , \147 , \363 );
mnand \mul_6_11_g6700/U$1 ( \435 , \433 , \434 );
mand \mul_6_11_g6612/U$3 ( \436 , \430 , \435 );
mand \mul_6_11_g6612/U$5 ( \437 , \424 , \429 );
mor \mul_6_11_g6612/U$2 ( \438 , \436 , \437 );
mxnor \mul_6_11_g6575/U$1 ( \439 , \423 , \438 );
mnot \mul_6_11_g6542/U$4 ( \440 , \439 );
mand \mul_6_11_g6542/U$2 ( \441 , \396 , \440 );
mand \mul_6_11_g6542/U$5 ( \442 , \439 , \395 );
mnor \mul_6_11_g6542/U$1 ( \443 , \441 , \442 );
mxor \mul_6_11_g6612/U$1 ( \444 , \424 , \429 );
mxor \mul_6_11_g6612/U$1_r1 ( \445 , \444 , \435 );
mnot \mul_6_11_g6611/U$1 ( \446 , \445 );
mnot \mul_6_11_g6571/U$3 ( \447 , \446 );
mxor \mul_6_11_g6618/U$4 ( \448 , \181 , \191 );
mand \mul_6_11_g6618/U$3 ( \449 , \448 , \200 );
mand \mul_6_11_g6618/U$5 ( \450 , \181 , \191 );
mor \mul_6_11_g6618/U$2 ( \451 , \449 , \450 );
mnot \fopt36720/U$1 ( \452 , \451 );
mnot \mul_6_11_g6571/U$4 ( \453 , \452 );
mor \mul_6_11_g6571/U$2 ( \454 , \447 , \453 );
mxor \mul_6_11_g6591/U$1 ( \455 , \378 , \384 );
mxor \mul_6_11_g6591/U$1_r1 ( \456 , \455 , \387 );
mnand \mul_6_11_g6571/U$1 ( \457 , \454 , \456 );
mnot \mul_6_11_g6920/U$2 ( \458 , \446 );
mnand \mul_6_11_g6920/U$1 ( \459 , \458 , \451 );
mnand \mul_6_11_g6559/U$1 ( \460 , \457 , \459 );
mnot \mul_6_11_g6553/U$1 ( \461 , \460 );
mnand \mul_6_11_g6514/U$1 ( \462 , \443 , \461 );
mxor \g36647/U$1 ( \463 , \445 , \452 );
mxor \g36647/U$1_r1 ( \464 , \463 , \456 );
mxor \mul_6_11_g6549/U$4 ( \465 , \170 , \174 );
mand \mul_6_11_g6549/U$3 ( \466 , \465 , \201 );
mand \mul_6_11_g6549/U$5 ( \467 , \170 , \174 );
mor \mul_6_11_g6549/U$2 ( \468 , \466 , \467 );
mnot \mul_6_11_g6548/U$1 ( \469 , \468 );
mnand \mul_6_11_g6533/U$1 ( \470 , \464 , \469 );
mand \mul_6_11_g6507/U$1 ( \471 , \462 , \470 );
mnot \mul_6_11_g6693/U$3 ( \472 , \374 );
mnot \mul_6_11_g6693/U$4 ( \473 , \359 );
mor \mul_6_11_g6693/U$2 ( \474 , \472 , \473 );
mxor \mul_6_11_g6847/U$1 ( \475 , \a[4] , \b[7] );
mnand \mul_6_11_g6744/U$1 ( \476 , \129 , \475 );
mnand \mul_6_11_g6693/U$1 ( \477 , \474 , \476 );
mnot \mul_6_11_g6687/U$3 ( \478 , \404 );
mnot \mul_6_11_g6687/U$4 ( \479 , \401 );
mor \mul_6_11_g6687/U$2 ( \480 , \478 , \479 );
mxor \mul_6_11_g6865/U$1 ( \481 , \a[2] , \b[9] );
mnand \mul_6_11_g6765/U$1 ( \482 , \400 , \481 );
mnand \mul_6_11_g6687/U$1 ( \483 , \480 , \482 );
mxor \mul_6_11_g6604/U$1 ( \484 , \477 , \483 );
mnot \mul_6_11_g6706/U$3 ( \485 , \367 );
mbuf \mul_6_11_g6762/U$1 ( \486 , \295 );
mnot \mul_6_11_g6706/U$4 ( \487 , \486 );
mor \mul_6_11_g6706/U$2 ( \488 , \485 , \487 );
mxor \mul_6_11_g6810/U$1 ( \489 , \a[8] , \b[3] );
mnand \mul_6_11_g6780/U$1 ( \490 , \147 , \489 );
mnand \mul_6_11_g6706/U$1 ( \491 , \488 , \490 );
mxor \mul_6_11_g6604/U$1_r1 ( \492 , \484 , \491 );
mnot \mul_6_11_g6572/U$3 ( \493 , \406 );
mnot \mul_6_11_g6572/U$4 ( \494 , \419 );
mor \mul_6_11_g6572/U$2 ( \495 , \493 , \494 );
mor \mul_6_11_g6579/U$2 ( \496 , \419 , \406 );
mnand \mul_6_11_g6579/U$1 ( \497 , \496 , \438 );
mnand \mul_6_11_g6572/U$1 ( \498 , \495 , \497 );
mxor \mul_6_11_g6525/U$1 ( \499 , \492 , \498 );
mand \mul_6_11_g6635/U$2 ( \500 , \412 , \418 );
mxor \mul_6_11_g6627/U$4 ( \501 , \354 , \361 );
mand \mul_6_11_g6627/U$3 ( \502 , \501 , \369 );
mand \mul_6_11_g6627/U$5 ( \503 , \354 , \361 );
mor \mul_6_11_g6627/U$2 ( \504 , \502 , \503 );
mxor \mul_6_11_g6565/U$1 ( \505 , \500 , \504 );
mxor \mul_6_11_g6836/U$1 ( \506 , \b[10] , \b[9] );
mand \mul_6_11_g6905/U$1 ( \507 , \506 , \a[0] );
mnot \mul_6_11_g6727/U$3 ( \508 , \352 );
mnot \mul_6_11_g6727/U$4 ( \509 , \120 );
mor \mul_6_11_g6727/U$2 ( \510 , \508 , \509 );
mxor \mul_6_11_g37182/U$1 ( \511 , \a[10] , \b[1] );
mnand \mul_6_11_g6774/U$1 ( \512 , \b[0] , \511 );
mnand \mul_6_11_g6727/U$1 ( \513 , \510 , \512 );
mxor \mul_6_11_g6605/U$1 ( \514 , \507 , \513 );
mnot \g37139/U$3 ( \515 , \195 );
mnot \g37139/U$4 ( \516 , \416 );
mor \g37139/U$2 ( \517 , \515 , \516 );
mxor \mul_6_11_g6830/U$1 ( \518 , \a[6] , \b[5] );
mnand \mul_6_11_g6712/U$1 ( \519 , \139 , \518 );
mnand \g37139/U$1 ( \520 , \517 , \519 );
mxor \mul_6_11_g6605/U$1_r1 ( \521 , \514 , \520 );
mxor \mul_6_11_g6565/U$1_r1 ( \522 , \505 , \521 );
mxnor \mul_6_11_g6525/U$1_r1 ( \523 , \499 , \522 );
mnot \mul_6_11_g6538/U$3 ( \524 , \393 );
mnot \mul_6_11_g6538/U$4 ( \525 , \439 );
mor \mul_6_11_g6538/U$2 ( \526 , \524 , \525 );
mbuf \fopt36721/U$1 ( \527 , \390 );
mnand \mul_6_11_g6538/U$1 ( \528 , \526 , \527 );
mor \mul_6_11_g6918/U$1 ( \529 , \439 , \393 );
mnand \mul_6_11_g6529/U$1 ( \530 , \528 , \529 );
mnot \fopt36739/U$1 ( \531 , \530 );
mnand \mul_6_11_g6511/U$1 ( \532 , \523 , \531 );
mnand \mul_6_11_g6499/U$1 ( \533 , \347 , \471 , \532 );
mnot \mul_6_11_g6509/U$3 ( \534 , \460 );
mnot \mul_6_11_g6523/U$1 ( \535 , \443 );
mnot \mul_6_11_g6509/U$4 ( \536 , \535 );
mor \mul_6_11_g6509/U$2 ( \537 , \534 , \536 );
mnot \mul_6_11_g6535/U$2 ( \538 , \469 );
mnot \mul_6_11_g6550/U$1 ( \539 , \464 );
mnand \mul_6_11_g6535/U$1 ( \540 , \538 , \539 );
mnand \mul_6_11_g6509/U$1 ( \541 , \537 , \540 );
mbuf \mul_6_11_g6513/U$1 ( \542 , \462 );
mnand \mul_6_11_g6501/U$1 ( \543 , \541 , \542 , \532 );
mnot \mul_6_11_g6912/U$2 ( \544 , \523 );
mnot \fopt36738/U$1 ( \545 , \531 );
mnand \mul_6_11_g6912/U$1 ( \546 , \544 , \545 );
mnand \mul_6_11_g6493/U$1 ( \547 , \533 , \543 , \546 );
mnand \mul_6_11_g6544/U$1 ( \548 , \522 , \492 );
mor \mul_6_11_g6537/U$2 ( \549 , \522 , \492 );
mnand \mul_6_11_g6537/U$1 ( \550 , \549 , \498 );
mnand \mul_6_11_g6527/U$1 ( \551 , \548 , \550 );
mxor \mul_6_11_g6605/U$4 ( \552 , \507 , \513 );
mand \mul_6_11_g6605/U$3 ( \553 , \552 , \520 );
mand \mul_6_11_g6605/U$5 ( \554 , \507 , \513 );
mor \mul_6_11_g6605/U$2 ( \555 , \553 , \554 );
mxor \mul_6_11_g6861/U$1 ( \556 , \b[11] , \b[10] );
mxor \mul_6_11_g6835/U$1 ( \557 , \a[0] , \b[11] );
mnand \mul_6_11_g6743/U$1 ( \558 , \556 , \557 );
mor \mul_6_11_g6678/U$2 ( \559 , \558 , \506 );
mxor \mul_6_11_g6853/U$1 ( \560 , \a[1] , \b[11] );
mnand \mul_6_11_g6761/U$1 ( \561 , \506 , \560 );
mnand \mul_6_11_g6678/U$1 ( \562 , \559 , \561 );
mor \mul_6_11_g6799/U$2 ( \563 , \a[0] , \b[10] );
mnand \mul_6_11_g6799/U$1 ( \564 , \563 , \b[9] );
mnand \mul_6_11_g6873/U$1 ( \565 , \a[0] , \b[10] );
mnand \mul_6_11_g6793/U$1 ( \566 , \564 , \565 , \b[11] );
mnot \mul_6_11_g6792/U$1 ( \567 , \566 );
mand \mul_6_11_g6651/U$2 ( \568 , \562 , \567 );
mnot \mul_6_11_g6651/U$4 ( \569 , \562 );
mand \mul_6_11_g6651/U$3 ( \570 , \569 , \566 );
mnor \mul_6_11_g6651/U$1 ( \571 , \568 , \570 );
mnot \mul_6_11_g6725/U$3 ( \572 , \511 );
mnot \mul_6_11_g6725/U$4 ( \573 , \120 );
mor \mul_6_11_g6725/U$2 ( \574 , \572 , \573 );
mxor \mul_6_11_g6823/U$1 ( \575 , \a[11] , \b[1] );
mnand \mul_6_11_g6771/U$1 ( \576 , \575 , \b[0] );
mnand \mul_6_11_g6725/U$1 ( \577 , \574 , \576 );
mnot \mul_6_11_g6724/U$1 ( \578 , \577 );
mand \mul_6_11_g6632/U$2 ( \579 , \571 , \578 );
mnot \mul_6_11_g6632/U$4 ( \580 , \571 );
mand \mul_6_11_g6632/U$3 ( \581 , \580 , \577 );
mnor \mul_6_11_g6632/U$1 ( \582 , \579 , \581 );
mxor \g37133/U$1 ( \583 , \555 , \582 );
mxor \mul_6_11_g6604/U$4 ( \584 , \477 , \483 );
mand \mul_6_11_g6604/U$3 ( \585 , \584 , \491 );
mand \mul_6_11_g6604/U$5 ( \586 , \477 , \483 );
mor \mul_6_11_g6604/U$2 ( \587 , \585 , \586 );
mxnor \g37133/U$1_r1 ( \588 , \583 , \587 );
mnot \mul_6_11_g6686/U$3 ( \589 , \481 );
mnot \mul_6_11_g6686/U$4 ( \590 , \401 );
mor \mul_6_11_g6686/U$2 ( \591 , \589 , \590 );
mxor \mul_6_11_g6864/U$1 ( \592 , \a[3] , \b[9] );
mnand \mul_6_11_g6766/U$1 ( \593 , \400 , \592 );
mnand \mul_6_11_g6686/U$1 ( \594 , \591 , \593 );
mnot \mul_6_11_g6668/U$3 ( \595 , \518 );
mnot \mul_6_11_g6668/U$4 ( \596 , \195 );
mor \mul_6_11_g6668/U$2 ( \597 , \595 , \596 );
mxor \mul_6_11_g6831/U$1 ( \598 , \a[7] , \b[5] );
mnand \mul_6_11_g6713/U$1 ( \599 , \139 , \598 );
mnand \mul_6_11_g6668/U$1 ( \600 , \597 , \599 );
mxnor \g36658/U$1 ( \601 , \594 , \600 );
mnot \mul_6_11_g6705/U$3 ( \602 , \489 );
mnot \mul_6_11_g6705/U$4 ( \603 , \486 );
mor \mul_6_11_g6705/U$2 ( \604 , \602 , \603 );
mnot \mul_6_11_g6878/U$2 ( \605 , \b[3] );
mnand \mul_6_11_g6878/U$1 ( \606 , \605 , \a[9] );
mnot \mul_6_11_g6781/U$3 ( \607 , \606 );
mnot \mul_6_11_g6872/U$2 ( \608 , \a[9] );
mnand \mul_6_11_g6872/U$1 ( \609 , \608 , \b[3] );
mnot \mul_6_11_g6781/U$4 ( \610 , \609 );
mor \mul_6_11_g6781/U$2 ( \611 , \607 , \610 );
mnand \mul_6_11_g6781/U$1 ( \612 , \611 , \147 );
mnand \mul_6_11_g6705/U$1 ( \613 , \604 , \612 );
mnot \mul_6_11_g6650/U$3 ( \614 , \613 );
mnot \mul_6_11_g6692/U$3 ( \615 , \475 );
mnot \mul_6_11_g6692/U$4 ( \616 , \374 );
mor \mul_6_11_g6692/U$2 ( \617 , \615 , \616 );
mxor \mul_6_11_g6848/U$1 ( \618 , \a[5] , \b[7] );
mnand \mul_6_11_g6745/U$1 ( \619 , \129 , \618 );
mnand \mul_6_11_g6692/U$1 ( \620 , \617 , \619 );
mnot \mul_6_11_g6691/U$1 ( \621 , \620 );
mnot \mul_6_11_g6650/U$4 ( \622 , \621 );
mand \mul_6_11_g6650/U$2 ( \623 , \614 , \622 );
mand \mul_6_11_g6650/U$5 ( \624 , \613 , \621 );
mnor \mul_6_11_g6650/U$1 ( \625 , \623 , \624 );
mnot \mul_6_11_g6929/U$2 ( \626 , \625 );
mxor \mul_6_11_g6929/U$1 ( \627 , \601 , \626 );
mnot \mul_6_11_g6607/U$1 ( \628 , \627 );
mand \mul_6_11_g6541/U$2 ( \629 , \588 , \628 );
mnot \mul_6_11_g6541/U$4 ( \630 , \588 );
mand \mul_6_11_g6541/U$3 ( \631 , \630 , \627 );
mnor \mul_6_11_g6541/U$1 ( \632 , \629 , \631 );
mxor \mul_6_11_g6565/U$4 ( \633 , \500 , \504 );
mand \mul_6_11_g6565/U$3 ( \634 , \633 , \521 );
mand \mul_6_11_g6565/U$5 ( \635 , \500 , \504 );
mor \mul_6_11_g6565/U$2 ( \636 , \634 , \635 );
mnot \mul_6_11_g6564/U$1 ( \637 , \636 );
mand \mul_6_11_g6521/U$2 ( \638 , \632 , \637 );
mnot \mul_6_11_g6521/U$4 ( \639 , \632 );
mand \mul_6_11_g6521/U$3 ( \640 , \639 , \636 );
mnor \mul_6_11_g6521/U$1 ( \641 , \638 , \640 );
mxor \mul_6_11_g36678/U$1 ( \642 , \551 , \641 );
mnot \mul_6_11_g6505/U$1 ( \643 , \642 );
mand \mul_6_11_g6489/U$2 ( \644 , \547 , \643 );
mnot \mul_6_11_g6489/U$4 ( \645 , \547 );
mand \mul_6_11_g6489/U$3 ( \646 , \645 , \642 );
mnor \mul_6_11_g6489/U$1 ( \647 , \644 , \646 );
mbuf \mul_6_11_g6488/U$1 ( \648 , \647 );
mbuf \g4836/U$1 ( \649 , \648 );
mnot \g4514/U$4 ( \650 , \649 );
mor \g4514/U$2 ( \651 , \99 , \650 );
mnot \mul_6_11_g6914/U$2 ( \652 , \535 );
mnor \mul_6_11_g6914/U$1 ( \653 , \652 , \461 );
mnot \mul_6_11_g6510/U$2 ( \654 , \653 );
mnand \mul_6_11_g6510/U$1 ( \655 , \654 , \542 );
mnot \mul_6_11_g6491/U$3 ( \656 , \655 );
mnot \mul_6_11_g6494/U$3 ( \657 , \470 );
mnot \mul_6_11_g6494/U$4 ( \658 , \347 );
mor \mul_6_11_g6494/U$2 ( \659 , \657 , \658 );
mnand \mul_6_11_g6536/U$1 ( \660 , \539 , \468 );
mbuf \fopt36958/U$1 ( \661 , \660 );
mnand \mul_6_11_g6494/U$1 ( \662 , \659 , \661 );
mnot \mul_6_11_g6491/U$4 ( \663 , \662 );
mor \mul_6_11_g6491/U$2 ( \664 , \656 , \663 );
mor \mul_6_11_g6491/U$5 ( \665 , \662 , \655 );
mnand \mul_6_11_g6491/U$1 ( \666 , \664 , \665 );
mbuf \g4798/U$1 ( \667 , \666 );
mand \g4523/U$2 ( \668 , \667 , \b[15] );
mnor \g36900/U$1 ( \669 , \a[11] , \d[11] );
mnot \g4597/U$2 ( \670 , \669 );
mnor \g4723/U$1 ( \671 , \a[8] , \a[7] , \a[6] , \a[5] );
mnor \g4744/U$1 ( \672 , \a[10] , \d[10] );
mnor \g4763/U$1 ( \673 , \a[9] , \d[9] );
mnor \g4752/U$1 ( \674 , \a[3] , \d[3] );
mnand \g4650/U$1 ( \675 , \671 , \672 , \673 , \674 );
mor \g4729/U$1 ( \676 , \a[15] , \a[4] , \d[8] , \d[7] );
mor \g4733/U$1 ( \677 , \d[6] , \d[5] , \d[15] , \d[4] );
mnor \g4628/U$1 ( \678 , \675 , \676 , \677 );
mand \g4654/U$2 ( \679 , \a[1] , \d[1] );
mnor \g4776/U$1 ( \680 , \a[1] , \d[1] );
mnor \g4770/U$1 ( \681 , \a[0] , \d[0] );
mnor \g4654/U$1 ( \682 , \679 , \680 , \681 );
mnor \g4765/U$1 ( \683 , \a[2] , \d[2] );
mnand \g37036/U$1 ( \684 , \a[0] , \d[0] );
mnand \g4603/U$1 ( \685 , \678 , \682 , \683 , \684 );
mor \g4760/U$1 ( \686 , \a[14] , \d[14] );
mnot \g4796/U$1 ( \687 , \d[12] );
mnot \g4843/U$1 ( \688 , \a[12] );
mnand \g4756/U$1 ( \689 , \687 , \688 );
mor \g4675/U$1 ( \690 , \686 , \689 , \d[13] );
mnor \g4597/U$1 ( \691 , \670 , \685 , \690 , \a[13] );
mnor \g4560/U$1 ( \692 , \691 , \d[15] );
mnot \g4532/U$3 ( \693 , \692 );
mnand \mul_6_11_g6916/U$1 ( \694 , \660 , \470 );
mxnor \g36646/U$1 ( \695 , \347 , \694 );
mnot \g4835/U$1 ( \696 , \695 );
mnot \g4834/U$1 ( \697 , \696 );
mnot \g4532/U$4 ( \698 , \697 );
mor \g4532/U$2 ( \699 , \693 , \698 );
mnot \mul_6_11_g6555/U$3 ( \700 , \262 );
mnot \mul_6_11_g6555/U$4 ( \701 , \266 );
mor \mul_6_11_g6555/U$2 ( \702 , \700 , \701 );
mnand \mul_6_11_g6555/U$1 ( \703 , \702 , \338 );
mbuf \mul_6_11_g6567/U$1 ( \704 , \335 );
mxnor \mul_6_11_g6917/U$1 ( \705 , \703 , \704 );
mnot \g4855/U$1 ( \706 , \705 );
mnot \g4854/U$1 ( \707 , \706 );
mnot \add_17_12_g6767/U$3 ( \708 , \b[15] );
mnot \add_17_12_g6767/U$4 ( \709 , \d[15] );
mand \add_17_12_g6767/U$2 ( \710 , \708 , \709 );
mand \add_17_12_g6767/U$5 ( \711 , \b[15] , \d[15] );
mnor \add_17_12_g6767/U$1 ( \712 , \710 , \711 );
mnot \add_17_12_g6684/U$3 ( \713 , \712 );
mnand \add_17_12_g6800/U$1 ( \714 , \b[0] , \d[0] );
mnand \add_17_12_g6777/U$1 ( \715 , \b[1] , \d[1] );
mnand \add_17_12_g6727/U$1 ( \716 , \714 , \715 );
mor \add_17_12_g6803/U$1 ( \717 , \b[1] , \d[1] );
mnor \add_17_12_g6784/U$1 ( \718 , \b[2] , \d[2] );
mnot \add_17_12_g6783/U$1 ( \719 , \718 );
mnand \add_17_12_g6725/U$1 ( \720 , \716 , \717 , \719 );
mnand \add_17_12_g6788/U$1 ( \721 , \b[3] , \d[3] );
mnand \add_17_12_g6778/U$1 ( \722 , \b[2] , \d[2] );
mnand \g37086/U$1 ( \723 , \720 , \721 , \722 );
mnot \g37085/U$3 ( \724 , \723 );
mnor \add_17_12_g6772/U$1 ( \725 , \b[5] , \d[5] );
mnor \add_17_12_g6797/U$1 ( \726 , \b[4] , \d[4] );
mnor \add_17_12_g6761/U$1 ( \727 , \725 , \726 );
mnor \add_17_12_g6770/U$1 ( \728 , \b[6] , \d[6] );
mnor \add_17_12_g6799/U$1 ( \729 , \b[7] , \d[7] );
mnor \add_17_12_g6765/U$1 ( \730 , \728 , \729 );
mnand \add_17_12_g6732/U$1 ( \731 , \727 , \730 );
mnor \add_17_12_g6786/U$1 ( \732 , \b[3] , \d[3] );
mnor \add_17_12_g6729/U$1 ( \733 , \731 , \732 );
mnot \g37085/U$4 ( \734 , \733 );
mor \g37085/U$2 ( \735 , \724 , \734 );
mnand \add_17_12_g6776/U$1 ( \736 , \b[7] , \d[7] );
mnot \add_17_12_g6722/U$3 ( \737 , \736 );
mnot \add_17_12_g6764/U$1 ( \738 , \730 );
mnot \add_17_12_g6722/U$4 ( \739 , \738 );
mor \add_17_12_g6722/U$2 ( \740 , \737 , \739 );
mnand \add_17_12_g6769/U$1 ( \741 , \b[6] , \d[6] );
mnand \add_17_12_g6785/U$1 ( \742 , \b[5] , \d[5] );
mnand \add_17_12_g6773/U$1 ( \743 , \b[4] , \d[4] );
mor \add_17_12_g6759/U$1 ( \744 , \725 , \743 );
mnand \g37087/U$1 ( \745 , \741 , \736 , \742 , \744 );
mnand \add_17_12_g6722/U$1 ( \746 , \740 , \745 );
mnand \g37085/U$1 ( \747 , \735 , \746 );
mnor \add_17_12_g6789/U$1 ( \748 , \b[11] , \d[11] );
mnor \add_17_12_g6780/U$1 ( \749 , \b[10] , \d[10] );
mnor \add_17_12_g6745/U$1 ( \750 , \748 , \749 );
mnor \add_17_12_g6791/U$1 ( \751 , \b[9] , \d[9] );
mnor \add_17_12_g6794/U$1 ( \752 , \b[8] , \d[8] );
mnor \add_17_12_g6752/U$1 ( \753 , \751 , \752 );
mand \add_17_12_g6735/U$1 ( \754 , \750 , \753 );
mnor \add_17_12_g6775/U$1 ( \755 , \b[14] , \d[14] );
mnot \add_17_12_g6734/U$2 ( \756 , \755 );
mnor \add_17_12_g6790/U$1 ( \757 , \b[13] , \d[13] );
mnor \add_17_12_g6795/U$1 ( \758 , \b[12] , \d[12] );
mnor \add_17_12_g6743/U$1 ( \759 , \757 , \758 );
mnand \add_17_12_g6734/U$1 ( \760 , \756 , \759 );
mnot \add_17_12_g6733/U$1 ( \761 , \760 );
mand \add_17_12_g6695/U$2 ( \762 , \747 , \754 , \761 );
mnand \add_17_12_g6793/U$1 ( \763 , \b[8] , \d[8] );
mor \add_17_12_g6738/U$2 ( \764 , \751 , \763 );
mnand \add_17_12_g6782/U$1 ( \765 , \b[9] , \d[9] );
mnand \add_17_12_g6738/U$1 ( \766 , \764 , \765 );
mnot \add_17_12_g6724/U$3 ( \767 , \766 );
mnot \add_17_12_g6724/U$4 ( \768 , \750 );
mor \add_17_12_g6724/U$2 ( \769 , \767 , \768 );
mnot \add_17_12_g6740/U$3 ( \770 , \748 );
mnand \add_17_12_g6774/U$1 ( \771 , \b[10] , \d[10] );
mnot \add_17_12_g6740/U$4 ( \772 , \771 );
mand \add_17_12_g6740/U$2 ( \773 , \770 , \772 );
mand \add_17_12_g6781/U$1 ( \774 , \b[11] , \d[11] );
mnor \add_17_12_g6740/U$1 ( \775 , \773 , \774 );
mnand \add_17_12_g6724/U$1 ( \776 , \769 , \775 );
mnot \add_17_12_g6723/U$1 ( \777 , \776 );
mor \add_17_12_g6715/U$2 ( \778 , \777 , \760 );
mnand \add_17_12_g6771/U$1 ( \779 , \b[12] , \d[12] );
mor \add_17_12_g6737/U$2 ( \780 , \757 , \779 );
mnand \add_17_12_g6792/U$1 ( \781 , \b[13] , \d[13] );
mnand \add_17_12_g6737/U$1 ( \782 , \780 , \781 );
mnot \add_17_12_g6736/U$1 ( \783 , \782 );
mor \add_17_12_g6715/U$3 ( \784 , \755 , \783 );
mnand \add_17_12_g6787/U$1 ( \785 , \b[14] , \d[14] );
mnand \add_17_12_g6715/U$1 ( \786 , \778 , \784 , \785 );
mnor \add_17_12_g6695/U$1 ( \787 , \762 , \786 );
mnot \add_17_12_g6684/U$4 ( \788 , \787 );
mor \add_17_12_g6684/U$2 ( \789 , \713 , \788 );
mor \add_17_12_g6684/U$5 ( \790 , \787 , \712 );
mnand \add_17_12_g6684/U$1 ( \791 , \789 , \790 );
mand \g4644/U$2 ( \792 , \707 , \791 );
mnot \add_16_12_g6767/U$3 ( \793 , \a[15] );
mnot \add_16_12_g6767/U$4 ( \794 , \c[15] );
mand \add_16_12_g6767/U$2 ( \795 , \793 , \794 );
mand \add_16_12_g6767/U$5 ( \796 , \a[15] , \c[15] );
mnor \add_16_12_g6767/U$1 ( \797 , \795 , \796 );
mnot \add_16_12_g6684/U$3 ( \798 , \797 );
mnand \add_16_12_g6800/U$1 ( \799 , \a[0] , \c[0] );
mnand \add_16_12_g6777/U$1 ( \800 , \a[1] , \c[1] );
mnand \add_16_12_g6727/U$1 ( \801 , \799 , \800 );
mor \add_16_12_g6803/U$1 ( \802 , \a[1] , \c[1] );
mnor \add_16_12_g6784/U$1 ( \803 , \a[2] , \c[2] );
mnot \add_16_12_g6783/U$1 ( \804 , \803 );
mnand \add_16_12_g6725/U$1 ( \805 , \801 , \802 , \804 );
mnand \add_16_12_g6788/U$1 ( \806 , \a[3] , \c[3] );
mnand \add_16_12_g6778/U$1 ( \807 , \a[2] , \c[2] );
mnand \g37089/U$1 ( \808 , \805 , \806 , \807 );
mnot \g37088/U$3 ( \809 , \808 );
mnor \add_16_12_g6772/U$1 ( \810 , \a[5] , \c[5] );
mnor \add_16_12_g6797/U$1 ( \811 , \a[4] , \c[4] );
mnor \add_16_12_g6761/U$1 ( \812 , \810 , \811 );
mnor \add_16_12_g6770/U$1 ( \813 , \a[6] , \c[6] );
mnor \add_16_12_g6799/U$1 ( \814 , \a[7] , \c[7] );
mnor \add_16_12_g6765/U$1 ( \815 , \813 , \814 );
mnand \add_16_12_g6732/U$1 ( \816 , \812 , \815 );
mnor \add_16_12_g6786/U$1 ( \817 , \a[3] , \c[3] );
mnor \add_16_12_g6729/U$1 ( \818 , \816 , \817 );
mnot \g37088/U$4 ( \819 , \818 );
mor \g37088/U$2 ( \820 , \809 , \819 );
mnand \add_16_12_g6776/U$1 ( \821 , \a[7] , \c[7] );
mnot \add_16_12_g6722/U$3 ( \822 , \821 );
mnot \add_16_12_g6764/U$1 ( \823 , \815 );
mnot \add_16_12_g6722/U$4 ( \824 , \823 );
mor \add_16_12_g6722/U$2 ( \825 , \822 , \824 );
mnand \add_16_12_g6769/U$1 ( \826 , \a[6] , \c[6] );
mnand \add_16_12_g6785/U$1 ( \827 , \a[5] , \c[5] );
mnand \add_16_12_g6773/U$1 ( \828 , \a[4] , \c[4] );
mor \add_16_12_g6759/U$1 ( \829 , \810 , \828 );
mnand \g37090/U$1 ( \830 , \826 , \821 , \827 , \829 );
mnand \add_16_12_g6722/U$1 ( \831 , \825 , \830 );
mnand \g37088/U$1 ( \832 , \820 , \831 );
mnor \add_16_12_g6789/U$1 ( \833 , \a[11] , \c[11] );
mnor \add_16_12_g6780/U$1 ( \834 , \a[10] , \c[10] );
mnor \add_16_12_g6745/U$1 ( \835 , \833 , \834 );
mnor \add_16_12_g6791/U$1 ( \836 , \a[9] , \c[9] );
mnor \add_16_12_g6794/U$1 ( \837 , \a[8] , \c[8] );
mnor \add_16_12_g6752/U$1 ( \838 , \836 , \837 );
mand \add_16_12_g6735/U$1 ( \839 , \835 , \838 );
mnor \add_16_12_g6775/U$1 ( \840 , \a[14] , \c[14] );
mnot \add_16_12_g6734/U$2 ( \841 , \840 );
mnor \add_16_12_g6790/U$1 ( \842 , \a[13] , \c[13] );
mnor \add_16_12_g6795/U$1 ( \843 , \a[12] , \c[12] );
mnor \add_16_12_g6743/U$1 ( \844 , \842 , \843 );
mnand \add_16_12_g6734/U$1 ( \845 , \841 , \844 );
mnot \add_16_12_g6733/U$1 ( \846 , \845 );
mand \add_16_12_g6695/U$2 ( \847 , \832 , \839 , \846 );
mnand \add_16_12_g6793/U$1 ( \848 , \a[8] , \c[8] );
mor \add_16_12_g6738/U$2 ( \849 , \836 , \848 );
mnand \add_16_12_g6782/U$1 ( \850 , \a[9] , \c[9] );
mnand \add_16_12_g6738/U$1 ( \851 , \849 , \850 );
mnot \add_16_12_g6724/U$3 ( \852 , \851 );
mnot \add_16_12_g6724/U$4 ( \853 , \835 );
mor \add_16_12_g6724/U$2 ( \854 , \852 , \853 );
mnot \add_16_12_g6740/U$3 ( \855 , \833 );
mnand \add_16_12_g6774/U$1 ( \856 , \a[10] , \c[10] );
mnot \add_16_12_g6740/U$4 ( \857 , \856 );
mand \add_16_12_g6740/U$2 ( \858 , \855 , \857 );
mand \add_16_12_g6781/U$1 ( \859 , \a[11] , \c[11] );
mnor \add_16_12_g6740/U$1 ( \860 , \858 , \859 );
mnand \add_16_12_g6724/U$1 ( \861 , \854 , \860 );
mnot \add_16_12_g6723/U$1 ( \862 , \861 );
mor \add_16_12_g6715/U$2 ( \863 , \862 , \845 );
mnand \add_16_12_g6771/U$1 ( \864 , \a[12] , \c[12] );
mor \add_16_12_g6737/U$2 ( \865 , \842 , \864 );
mnand \add_16_12_g6792/U$1 ( \866 , \a[13] , \c[13] );
mnand \add_16_12_g6737/U$1 ( \867 , \865 , \866 );
mnot \add_16_12_g6736/U$1 ( \868 , \867 );
mor \add_16_12_g6715/U$3 ( \869 , \840 , \868 );
mnand \add_16_12_g6787/U$1 ( \870 , \a[14] , \c[14] );
mnand \add_16_12_g6715/U$1 ( \871 , \863 , \869 , \870 );
mnor \add_16_12_g6695/U$1 ( \872 , \847 , \871 );
mnot \add_16_12_g6684/U$4 ( \873 , \872 );
mor \add_16_12_g6684/U$2 ( \874 , \798 , \873 );
mor \add_16_12_g6684/U$5 ( \875 , \872 , \797 );
mnand \add_16_12_g6684/U$1 ( \876 , \874 , \875 );
mnot \g4670/U$3 ( \877 , \876 );
mnand \mul_6_11_g6586/U$1 ( \878 , \334 , \291 );
mxnor \mul_6_11_g6574/U$1 ( \879 , \878 , \329 );
mbuf \g4841/U$1 ( \880 , \879 );
mnot \g4670/U$4 ( \881 , \880 );
mor \g4670/U$2 ( \882 , \877 , \881 );
mor \mul_6_11_g6720/U$2 ( \883 , \314 , \208 );
mnand \mul_6_11_g6720/U$1 ( \884 , \883 , \318 );
mand \mul_6_11_g6904/U$1 ( \885 , \320 , \884 );
mnot \g4794/U$1 ( \886 , \885 );
mnot \g4711/U$3 ( \887 , \886 );
mnot \g4795/U$1 ( \888 , \b[15] );
mnot \g4711/U$4 ( \889 , \888 );
mand \g4711/U$2 ( \890 , \887 , \889 );
mnand \mul_6_11_g6628/U$1 ( \891 , \328 , \302 );
mxnor \mul_6_11_g6921/U$1 ( \892 , \891 , \324 );
mnot \g4828/U$1 ( \893 , \892 );
mnot \g4827/U$1 ( \894 , \893 );
mand \g4711/U$5 ( \895 , \894 , \d[15] );
mnor \g4711/U$1 ( \896 , \890 , \895 );
mnand \g4670/U$1 ( \897 , \882 , \896 );
mnor \g4644/U$1 ( \898 , \792 , \897 );
mnand \g4532/U$1 ( \899 , \699 , \898 );
mnor \g4523/U$1 ( \900 , \668 , \899 );
mnand \g4514/U$1 ( \901 , \651 , \900 );
mnot \g4602/U$1 ( \902 , \685 );
mbuf \g4832/U$1 ( \903 , \697 );
mand \g4573/U$2 ( \904 , \902 , \903 );
mnot \mul_6_11_g6662/U$2 ( \905 , \312 );
mnand \mul_6_11_g6662/U$1 ( \906 , \905 , \323 );
mxor \mul_6_11_g6927/U$1 ( \907 , \906 , \320 );
mnot \g4885/U$1 ( \908 , \907 );
mnot \g4884/U$1 ( \909 , \908 );
mnor \g4573/U$1 ( \910 , \904 , \909 );
mnot \g36779/U$3 ( \911 , \471 );
mnot \g36779/U$4 ( \912 , \347 );
mor \g36779/U$2 ( \913 , \911 , \912 );
mnand \mul_6_11_g6504/U$1 ( \914 , \541 , \542 );
mnand \g36779/U$1 ( \915 , \913 , \914 );
mxnor \g36833/U$1 ( \916 , \523 , \531 );
mnot \mul_6_11_g36945/U$1 ( \917 , \916 );
mand \g36944/U$2 ( \918 , \915 , \917 );
mnot \g36944/U$4 ( \919 , \915 );
mand \g36944/U$3 ( \920 , \919 , \916 );
mnor \g36944/U$1 ( \921 , \918 , \920 );
mbuf \g4858/U$1 ( \922 , \921 );
mnand \g4785/U$1 ( \923 , \922 , \b[15] );
mand \g4530/U$2 ( \924 , \910 , \923 );
mnot \g4867/U$1 ( \925 , \c[15] );
mnor \g4530/U$1 ( \926 , \924 , \925 );
mnor \g4512/U$1 ( \927 , \901 , \926 );
mxor \g36634/U$1 ( \928 , \d[5] , \a[6] );
mnot \mul_18_12_g22638/U$3 ( \929 , \928 );
mxor \mul_18_12_g22870/U$1 ( \930 , \d[5] , \d[4] );
mnot \mul_18_12_g22722/U$2 ( \931 , \930 );
mxor \mul_18_12_g36670/U$1 ( \932 , \d[4] , \d[3] );
mnor \mul_18_12_g22722/U$1 ( \933 , \931 , \932 );
mnot \mul_18_12_g22638/U$4 ( \934 , \933 );
mor \mul_18_12_g22638/U$2 ( \935 , \929 , \934 );
mbuf \mul_18_12_g22851/U$1 ( \936 , \932 );
mxor \g36633/U$1 ( \937 , \d[5] , \a[7] );
mnand \mul_18_12_g22710/U$1 ( \938 , \936 , \937 );
mnand \mul_18_12_g22638/U$1 ( \939 , \935 , \938 );
mxor \mul_18_12_g22930/U$1 ( \940 , \a[0] , \d[11] );
mnot \mul_18_12_g22615/U$3 ( \941 , \940 );
mxnor \mul_18_12_g36668/U$1 ( \942 , \d[11] , \d[10] );
mxor \mul_18_12_g22875/U$1 ( \943 , \d[10] , \d[9] );
mnor \mul_18_12_g22811/U$1 ( \944 , \942 , \943 );
mnot \mul_18_12_g22615/U$4 ( \945 , \944 );
mor \mul_18_12_g22615/U$2 ( \946 , \941 , \945 );
mxor \mul_18_12_g22876/U$1 ( \947 , \d[10] , \d[9] );
mxor \mul_18_12_g22944/U$1 ( \948 , \a[1] , \d[11] );
mnand \mul_18_12_g22711/U$1 ( \949 , \947 , \948 );
mnand \mul_18_12_g22615/U$1 ( \950 , \946 , \949 );
mnot \mul_18_12_g22614/U$1 ( \951 , \950 );
mxor \g36622/U$1 ( \952 , \939 , \951 );
mor \mul_18_12_g22818/U$2 ( \953 , \a[0] , \d[10] );
mnand \mul_18_12_g22818/U$1 ( \954 , \953 , \d[9] );
mnand \mul_18_12_g22956/U$1 ( \955 , \a[0] , \d[10] );
mand \mul_18_12_g23029/U$1 ( \956 , \954 , \955 , \d[11] );
mxor \mul_18_12_g22883/U$1 ( \957 , \a[8] , \d[3] );
mnot \mul_18_12_g22662/U$3 ( \958 , \957 );
mxor \mul_18_12_g23018/U$1 ( \959 , \d[2] , \d[1] );
mnot \fopt36726/U$1 ( \960 , \959 );
mxor \g36747/U$1 ( \961 , \d[3] , \d[2] );
mand \mul_18_12_g22761/U$1 ( \962 , \960 , \961 );
mnot \mul_18_12_g22662/U$4 ( \963 , \962 );
mor \mul_18_12_g22662/U$2 ( \964 , \958 , \963 );
mbuf \fopt36728/U$1 ( \965 , \959 );
mxor \mul_18_12_g22882/U$1 ( \966 , \a[9] , \d[3] );
mnand \mul_18_12_g22729/U$1 ( \967 , \965 , \966 );
mnand \mul_18_12_g22662/U$1 ( \968 , \964 , \967 );
mxor \mul_18_12_g22527/U$1 ( \969 , \956 , \968 );
mxnor \g36622/U$1_r1 ( \970 , \952 , \969 );
mor \mul_18_12_g22819/U$2 ( \971 , \a[0] , \d[8] );
mnand \mul_18_12_g22819/U$1 ( \972 , \971 , \d[7] );
mnand \mul_18_12_g22951/U$1 ( \973 , \a[0] , \d[8] );
mnand \mul_18_12_g22799/U$1 ( \974 , \972 , \973 , \d[9] );
mnot \mul_18_12_g23072/U$2 ( \975 , \974 );
mxor \mul_18_12_g22895/U$1 ( \976 , \a[6] , \d[3] );
mnot \mul_18_12_g22666/U$3 ( \977 , \976 );
mxor \mul_18_12_g36748/U$1 ( \978 , \d[3] , \d[2] );
mnot \mul_18_12_g22760/U$2 ( \979 , \978 );
mnor \mul_18_12_g22760/U$1 ( \980 , \979 , \959 );
mnot \mul_18_12_g22666/U$4 ( \981 , \980 );
mor \mul_18_12_g22666/U$2 ( \982 , \977 , \981 );
mxor \mul_18_12_g22893/U$1 ( \983 , \a[7] , \d[3] );
mnand \mul_18_12_g22732/U$1 ( \984 , \965 , \983 );
mnand \mul_18_12_g22666/U$1 ( \985 , \982 , \984 );
mnand \mul_18_12_g23072/U$1 ( \986 , \975 , \985 );
mnot \mul_18_12_g22416/U$3 ( \987 , \986 );
mnand \mul_18_12_g36751/U$1 ( \988 , \943 , \a[0] );
mnot \mul_18_12_g22776/U$1 ( \989 , \988 );
mnand \mul_18_12_g22716/U$1 ( \990 , \983 , \978 );
mor \g37125/U$2 ( \991 , \959 , \990 );
mnand \mul_18_12_g22731/U$1 ( \992 , \959 , \957 );
mnand \g37125/U$1 ( \993 , \991 , \992 );
mxor \mul_18_12_g22475/U$1 ( \994 , \989 , \993 );
mxor \g36640/U$1 ( \995 , \d[7] , \a[3] );
mnot \mul_18_12_g22626/U$3 ( \996 , \995 );
mxnor \mul_18_12_g23032/U$1 ( \997 , \d[7] , \d[6] );
mxor \mul_18_12_g36669/U$1 ( \998 , \d[6] , \d[5] );
mnor \mul_18_12_g22707/U$1 ( \999 , \997 , \998 );
mnot \mul_18_12_g22626/U$4 ( \1000 , \999 );
mor \mul_18_12_g22626/U$2 ( \1001 , \996 , \1000 );
mnot \mul_18_12_g22868/U$1 ( \1002 , \998 );
mnot \mul_18_12_g22864/U$1 ( \1003 , \1002 );
mxor \g36635/U$1 ( \1004 , \d[7] , \a[4] );
mnand \mul_18_12_g22705/U$1 ( \1005 , \1003 , \1004 );
mnand \mul_18_12_g22626/U$1 ( \1006 , \1001 , \1005 );
mxnor \mul_18_12_g22475/U$1_r1 ( \1007 , \994 , \1006 );
mnot \mul_18_12_g22416/U$4 ( \1008 , \1007 );
mor \mul_18_12_g22416/U$2 ( \1009 , \987 , \1008 );
mnot \mul_18_12_g23019/U$2 ( \1010 , \d[0] );
mnand \mul_18_12_g23019/U$1 ( \1011 , \1010 , \d[1] );
mnot \fopt36813/U$1 ( \1012 , \1011 );
mxor \g36629/U$1 ( \1013 , \d[1] , \a[8] );
mand \g37283/U$2 ( \1014 , \1012 , \1013 );
mxor \g36630/U$1 ( \1015 , \d[1] , \a[9] );
mand \g37283/U$3 ( \1016 , \1015 , \d[0] );
mnor \g37283/U$1 ( \1017 , \1014 , \1016 );
mnot \mul_18_12_g22698/U$1 ( \1018 , \1017 );
mnot \mul_18_12_g22499/U$3 ( \1019 , \1018 );
mxor \g36642/U$1 ( \1020 , \d[9] , \a[0] );
mnot \mul_18_12_g22573/U$3 ( \1021 , \1020 );
mor \mul_18_12_g23034/U$1 ( \1022 , \d[9] , \d[8] );
mnot \mul_18_12_g23011/U$2 ( \1023 , \d[7] );
mnand \mul_18_12_g23011/U$1 ( \1024 , \1023 , \d[8] );
mnand \mul_18_12_g37175/U$1 ( \1025 , \d[9] , \d[7] );
mand \mul_18_12_g22678/U$1 ( \1026 , \1022 , \1024 , \1025 );
mnot \mul_18_12_g22573/U$4 ( \1027 , \1026 );
mor \mul_18_12_g22573/U$2 ( \1028 , \1021 , \1027 );
mxor \mul_18_12_g22823/U$1 ( \1029 , \d[8] , \d[7] );
mxor \g36643/U$1 ( \1030 , \d[9] , \a[1] );
mnand \mul_18_12_g22670/U$1 ( \1031 , \1029 , \1030 );
mnand \mul_18_12_g22573/U$1 ( \1032 , \1028 , \1031 );
mnot \mul_18_12_g22499/U$4 ( \1033 , \1032 );
mor \mul_18_12_g22499/U$2 ( \1034 , \1019 , \1033 );
mor \mul_18_12_g22520/U$2 ( \1035 , \1032 , \1018 );
mxor \g36639/U$1 ( \1036 , \d[7] , \a[2] );
mnot \mul_18_12_g22622/U$3 ( \1037 , \1036 );
mnor \mul_18_12_g22706/U$1 ( \1038 , \997 , \998 );
mnot \mul_18_12_g22622/U$4 ( \1039 , \1038 );
mor \mul_18_12_g22622/U$2 ( \1040 , \1037 , \1039 );
mnot \mul_18_12_g23074/U$2 ( \1041 , \1002 );
mnand \mul_18_12_g23074/U$1 ( \1042 , \1041 , \995 );
mnand \mul_18_12_g22622/U$1 ( \1043 , \1040 , \1042 );
mnand \mul_18_12_g22520/U$1 ( \1044 , \1035 , \1043 );
mnand \mul_18_12_g22499/U$1 ( \1045 , \1034 , \1044 );
mnand \mul_18_12_g22416/U$1 ( \1046 , \1009 , \1045 );
mnot \mul_18_12_g23055/U$2 ( \1047 , \986 );
mnot \mul_18_12_g22466/U$1 ( \1048 , \1007 );
mnand \mul_18_12_g23055/U$1 ( \1049 , \1047 , \1048 );
mnand \mul_18_12_g22408/U$1 ( \1050 , \1046 , \1049 );
mxor \mul_18_12_g23046/U$1 ( \1051 , \970 , \1050 );
mxor \mul_18_12_g22935/U$1 ( \1052 , \a[2] , \d[9] );
mnot \mul_18_12_g22571/U$3 ( \1053 , \1052 );
mnot \mul_18_12_g22824/U$3 ( \1054 , \d[7] );
mnot \mul_18_12_g23015/U$1 ( \1055 , \d[8] );
mnot \mul_18_12_g22824/U$4 ( \1056 , \1055 );
mor \mul_18_12_g22824/U$2 ( \1057 , \1054 , \1056 );
mnand \mul_18_12_g22824/U$1 ( \1058 , \1057 , \1024 );
mnot \mul_18_12_g22571/U$4 ( \1059 , \1058 );
mor \mul_18_12_g22571/U$2 ( \1060 , \1053 , \1059 );
mnand \mul_18_12_g36834/U$1 ( \1061 , \1026 , \1030 );
mnand \mul_18_12_g22571/U$1 ( \1062 , \1060 , \1061 );
mnot \g37121/U$3 ( \1063 , \1062 );
mnot \mul_18_12_g22695/U$3 ( \1064 , \1015 );
mnot \fopt36810/U$1 ( \1065 , \1011 );
mnot \mul_18_12_g22695/U$4 ( \1066 , \1065 );
mor \mul_18_12_g22695/U$2 ( \1067 , \1064 , \1066 );
mxor \mul_18_12_g22845/U$1 ( \1068 , \a[10] , \d[1] );
mnand \mul_18_12_g22749/U$1 ( \1069 , \1068 , \d[0] );
mnand \mul_18_12_g22695/U$1 ( \1070 , \1067 , \1069 );
mnot \g37121/U$4 ( \1071 , \1070 );
mor \g37121/U$2 ( \1072 , \1063 , \1071 );
mor \mul_18_12_g22470/U$2 ( \1073 , \1070 , \1062 );
mxor \mul_18_12_g22910/U$1 ( \1074 , \a[5] , \d[5] );
mnot \mul_18_12_g22652/U$3 ( \1075 , \1074 );
mnot \mul_18_12_g22652/U$4 ( \1076 , \933 );
mor \mul_18_12_g22652/U$2 ( \1077 , \1075 , \1076 );
mnand \mul_18_12_g22763/U$1 ( \1078 , \936 , \928 );
mnand \mul_18_12_g22652/U$1 ( \1079 , \1077 , \1078 );
mnand \mul_18_12_g22470/U$1 ( \1080 , \1073 , \1079 );
mnand \g37121/U$1 ( \1081 , \1072 , \1080 );
mnot \g37166/U$2 ( \1082 , \993 );
mnand \g37166/U$1 ( \1083 , \1082 , \988 );
mnot \g37165/U$3 ( \1084 , \1083 );
mnot \g37165/U$4 ( \1085 , \1006 );
mor \g37165/U$2 ( \1086 , \1084 , \1085 );
mnand \mul_18_12_g22553/U$1 ( \1087 , \993 , \989 );
mnand \g37165/U$1 ( \1088 , \1086 , \1087 );
mxor \g36645/U$1 ( \1089 , \1081 , \1088 );
mnot \mul_18_12_g22684/U$3 ( \1090 , \1068 );
mnot \mul_18_12_g22684/U$4 ( \1091 , \1065 );
mor \mul_18_12_g22684/U$2 ( \1092 , \1090 , \1091 );
mxor \mul_18_12_g22844/U$1 ( \1093 , \a[11] , \d[1] );
mnand \mul_18_12_g22738/U$1 ( \1094 , \1093 , \d[0] );
mnand \mul_18_12_g22684/U$1 ( \1095 , \1092 , \1094 );
mnot \mul_18_12_g22683/U$1 ( \1096 , \1095 );
mnot \mul_18_12_g22536/U$3 ( \1097 , \1096 );
mnot \mul_18_12_g22630/U$3 ( \1098 , \1004 );
mnot \mul_18_12_g22630/U$4 ( \1099 , \1038 );
mor \mul_18_12_g22630/U$2 ( \1100 , \1098 , \1099 );
mxor \mul_18_12_g22911/U$1 ( \1101 , \a[5] , \d[7] );
mnand \mul_18_12_g22745/U$1 ( \1102 , \1003 , \1101 );
mnand \mul_18_12_g22630/U$1 ( \1103 , \1100 , \1102 );
mnot \mul_18_12_g22536/U$4 ( \1104 , \1103 );
mor \mul_18_12_g22536/U$2 ( \1105 , \1097 , \1104 );
mnot \mul_18_12_g22552/U$2 ( \1106 , \1103 );
mnand \mul_18_12_g22552/U$1 ( \1107 , \1106 , \1095 );
mnand \mul_18_12_g22536/U$1 ( \1108 , \1105 , \1107 );
mand \g37127/U$1 ( \1109 , \1024 , \1022 , \1025 );
mnot \mul_18_12_g22677/U$1 ( \1110 , \1109 );
mnot \mul_18_12_g22564/U$3 ( \1111 , \1110 );
mnot \mul_18_12_g22934/U$1 ( \1112 , \1052 );
mnot \mul_18_12_g22564/U$4 ( \1113 , \1112 );
mand \mul_18_12_g22564/U$2 ( \1114 , \1111 , \1113 );
mxor \mul_18_12_g22936/U$1 ( \1115 , \a[3] , \d[9] );
mand \mul_18_12_g22564/U$5 ( \1116 , \1058 , \1115 );
mnor \mul_18_12_g22564/U$1 ( \1117 , \1114 , \1116 );
mnot \fopt36709/U$1 ( \1118 , \1117 );
mbuf \fopt36708/U$1 ( \1119 , \1118 );
mand \mul_18_12_g22509/U$2 ( \1120 , \1108 , \1119 );
mnot \mul_18_12_g22509/U$4 ( \1121 , \1108 );
mnot \fopt36707/U$1 ( \1122 , \1119 );
mand \mul_18_12_g22509/U$3 ( \1123 , \1121 , \1122 );
mnor \mul_18_12_g22509/U$1 ( \1124 , \1120 , \1123 );
mxnor \g36645/U$1_r1 ( \1125 , \1089 , \1124 );
mxor \mul_18_12_g23046/U$1_r1 ( \1126 , \1051 , \1125 );
mxor \g37131/U$1 ( \1127 , \1062 , \1070 );
mxnor \g37131/U$1_r1 ( \1128 , \1127 , \1079 );
mxor \mul_18_12_g22908/U$1 ( \1129 , \a[4] , \d[5] );
mand \g37072/U$2 ( \1130 , \933 , \1129 );
mand \mul_18_12_g23075/U$1 ( \1131 , \936 , \1074 );
mnor \g37072/U$1 ( \1132 , \1130 , \1131 );
mnot \mul_18_12_g22534/U$3 ( \1133 , \985 );
mnot \mul_18_12_g22534/U$4 ( \1134 , \974 );
mand \mul_18_12_g22534/U$2 ( \1135 , \1133 , \1134 );
mand \mul_18_12_g22534/U$5 ( \1136 , \985 , \974 );
mnor \mul_18_12_g22534/U$1 ( \1137 , \1135 , \1136 );
mxor \mul_18_12_g22393/U$4 ( \1138 , \1132 , \1137 );
mnand \mul_18_12_g22675/U$1 ( \1139 , \1029 , \a[0] );
mxor \g36631/U$1 ( \1140 , \d[1] , \a[7] );
mand \g37128/U$2 ( \1141 , \1012 , \1140 );
mand \g37128/U$3 ( \1142 , \1013 , \d[0] );
mnor \g37128/U$1 ( \1143 , \1141 , \1142 );
mxor \mul_18_12_g22489/U$4 ( \1144 , \1139 , \1143 );
mxor \mul_18_12_g22937/U$1 ( \1145 , \a[1] , \d[7] );
mand \mul_18_12_g22623/U$2 ( \1146 , \1038 , \1145 );
mand \mul_18_12_g22623/U$3 ( \1147 , \1003 , \1036 );
mnor \mul_18_12_g22623/U$1 ( \1148 , \1146 , \1147 );
mand \mul_18_12_g22489/U$3 ( \1149 , \1144 , \1148 );
mand \mul_18_12_g22489/U$5 ( \1150 , \1139 , \1143 );
mor \mul_18_12_g22489/U$2 ( \1151 , \1149 , \1150 );
mand \mul_18_12_g22393/U$3 ( \1152 , \1138 , \1151 );
mand \mul_18_12_g22393/U$5 ( \1153 , \1132 , \1137 );
mor \mul_18_12_g22393/U$2 ( \1154 , \1152 , \1153 );
mxor \mul_18_12_g22328/U$4 ( \1155 , \1128 , \1154 );
mxor \mul_18_12_g22409/U$1 ( \1156 , \986 , \1045 );
mxor \mul_18_12_g22409/U$1_r1 ( \1157 , \1156 , \1048 );
mand \mul_18_12_g22328/U$3 ( \1158 , \1155 , \1157 );
mand \mul_18_12_g22328/U$5 ( \1159 , \1128 , \1154 );
mor \mul_18_12_g22328/U$2 ( \1160 , \1158 , \1159 );
mnand \mul_18_12_g22287/U$1 ( \1161 , \1126 , \1160 );
mxor \mul_18_12_g22328/U$1 ( \1162 , \1128 , \1154 );
mxor \mul_18_12_g22328/U$1_r1 ( \1163 , \1162 , \1157 );
mnot \mul_18_12_g22535/U$3 ( \1164 , \1017 );
mnot \mul_18_12_g22535/U$4 ( \1165 , \1043 );
mor \mul_18_12_g22535/U$2 ( \1166 , \1164 , \1165 );
mnot \mul_18_12_g22551/U$2 ( \1167 , \1043 );
mnand \mul_18_12_g22551/U$1 ( \1168 , \1167 , \1018 );
mnand \mul_18_12_g22535/U$1 ( \1169 , \1166 , \1168 );
mxor \mul_18_12_g23058/U$1 ( \1170 , \1169 , \1032 );
mnot \mul_18_12_g23052/U$2 ( \1171 , \1170 );
mnot \mul_18_12_g22686/U$3 ( \1172 , \1012 );
mxor \g36632/U$1 ( \1173 , \d[1] , \a[6] );
mnot \mul_18_12_g22686/U$4 ( \1174 , \1173 );
mor \mul_18_12_g22686/U$2 ( \1175 , \1172 , \1174 );
mnand \mul_18_12_g22717/U$1 ( \1176 , \1140 , \d[0] );
mnand \mul_18_12_g22686/U$1 ( \1177 , \1175 , \1176 );
mor \mul_18_12_g22820/U$2 ( \1178 , \a[0] , \d[6] );
mnand \mul_18_12_g22820/U$1 ( \1179 , \1178 , \d[5] );
mnand \mul_18_12_g22954/U$1 ( \1180 , \a[0] , \d[6] );
mand \mul_18_12_g22797/U$1 ( \1181 , \1179 , \1180 , \d[7] );
mnand \mul_18_12_g22592/U$1 ( \1182 , \1177 , \1181 );
mxor \mul_18_12_g22919/U$1 ( \1183 , \a[3] , \d[5] );
mnot \mul_18_12_g22642/U$3 ( \1184 , \1183 );
mnot \mul_18_12_g22723/U$2 ( \1185 , \930 );
mnor \mul_18_12_g22723/U$1 ( \1186 , \1185 , \932 );
mnot \mul_18_12_g22642/U$4 ( \1187 , \1186 );
mor \mul_18_12_g22642/U$2 ( \1188 , \1184 , \1187 );
mnand \mul_18_12_g22718/U$1 ( \1189 , \936 , \1129 );
mnand \mul_18_12_g22642/U$1 ( \1190 , \1188 , \1189 );
mnot \mul_18_12_g22641/U$1 ( \1191 , \1190 );
mnand \mul_18_12_g22513/U$1 ( \1192 , \1182 , \1191 );
mxor \mul_18_12_g22903/U$1 ( \1193 , \a[5] , \d[3] );
mnot \mul_18_12_g22659/U$3 ( \1194 , \1193 );
mnot \mul_18_12_g22659/U$4 ( \1195 , \962 );
mor \mul_18_12_g22659/U$2 ( \1196 , \1194 , \1195 );
mnand \mul_18_12_g22724/U$1 ( \1197 , \965 , \976 );
mnand \mul_18_12_g22659/U$1 ( \1198 , \1196 , \1197 );
mand \mul_18_12_g22441/U$2 ( \1199 , \1192 , \1198 );
mnot \mul_18_12_g22544/U$1 ( \1200 , \1182 );
mand \g37046/U$1 ( \1201 , \1200 , \1190 );
mnor \mul_18_12_g22441/U$1 ( \1202 , \1199 , \1201 );
mnand \mul_18_12_g23052/U$1 ( \1203 , \1171 , \1202 );
mnot \mul_18_12_g22341/U$3 ( \1204 , \1203 );
mxor \mul_18_12_g22393/U$1 ( \1205 , \1132 , \1137 );
mxor \mul_18_12_g22393/U$1_r1 ( \1206 , \1205 , \1151 );
mnot \mul_18_12_g22392/U$1 ( \1207 , \1206 );
mnot \mul_18_12_g22341/U$4 ( \1208 , \1207 );
mor \mul_18_12_g22341/U$2 ( \1209 , \1204 , \1208 );
mnot \mul_18_12_g23048/U$2 ( \1210 , \1202 );
mnand \mul_18_12_g23048/U$1 ( \1211 , \1210 , \1170 );
mnand \mul_18_12_g22341/U$1 ( \1212 , \1209 , \1211 );
mnot \mul_18_12_g22334/U$1 ( \1213 , \1212 );
mnand \mul_18_12_g22314/U$1 ( \1214 , \1163 , \1213 );
mxor \mul_18_12_g22489/U$1 ( \1215 , \1139 , \1143 );
mxor \mul_18_12_g22489/U$1_r1 ( \1216 , \1215 , \1148 );
mnot \mul_18_12_g22486/U$1 ( \1217 , \1216 );
mnot \mul_18_12_g22429/U$3 ( \1218 , \1217 );
mxor \mul_18_12_g22904/U$1 ( \1219 , \a[4] , \d[3] );
mnot \mul_18_12_g22664/U$3 ( \1220 , \1219 );
mnot \mul_18_12_g22664/U$4 ( \1221 , \962 );
mor \mul_18_12_g22664/U$2 ( \1222 , \1220 , \1221 );
mnand \mul_18_12_g22742/U$1 ( \1223 , \965 , \1193 );
mnand \mul_18_12_g22664/U$1 ( \1224 , \1222 , \1223 );
mxor \mul_18_12_g22920/U$1 ( \1225 , \a[2] , \d[5] );
mnot \mul_18_12_g22648/U$3 ( \1226 , \1225 );
mnot \mul_18_12_g22648/U$4 ( \1227 , \1186 );
mor \mul_18_12_g22648/U$2 ( \1228 , \1226 , \1227 );
mnand \mul_18_12_g22756/U$1 ( \1229 , \936 , \1183 );
mnand \mul_18_12_g22648/U$1 ( \1230 , \1228 , \1229 );
mor \mul_18_12_g22494/U$2 ( \1231 , \1224 , \1230 );
mxor \mul_18_12_g22943/U$1 ( \1232 , \a[0] , \d[7] );
mnot \mul_18_12_g22628/U$3 ( \1233 , \1232 );
mnot \mul_18_12_g22628/U$4 ( \1234 , \999 );
mor \mul_18_12_g22628/U$2 ( \1235 , \1233 , \1234 );
mnand \mul_18_12_g22725/U$1 ( \1236 , \1003 , \1145 );
mnand \mul_18_12_g22628/U$1 ( \1237 , \1235 , \1236 );
mnand \mul_18_12_g22494/U$1 ( \1238 , \1231 , \1237 );
mnand \mul_18_12_g22556/U$1 ( \1239 , \1224 , \1230 );
mnand \mul_18_12_g22473/U$1 ( \1240 , \1238 , \1239 );
mnot \mul_18_12_g22456/U$1 ( \1241 , \1240 );
mnot \mul_18_12_g22429/U$4 ( \1242 , \1241 );
mor \mul_18_12_g22429/U$2 ( \1243 , \1218 , \1242 );
mnand \mul_18_12_g22431/U$1 ( \1244 , \1240 , \1216 );
mnand \mul_18_12_g22429/U$1 ( \1245 , \1243 , \1244 );
mnot \mul_18_12_g22504/U$3 ( \1246 , \1191 );
mnot \mul_18_12_g22504/U$4 ( \1247 , \1200 );
mor \mul_18_12_g22504/U$2 ( \1248 , \1246 , \1247 );
mor \mul_18_12_g22504/U$5 ( \1249 , \1200 , \1191 );
mnand \mul_18_12_g22504/U$1 ( \1250 , \1248 , \1249 );
mnot \fopt36706/U$1 ( \1251 , \1198 );
mand \mul_18_12_g22442/U$2 ( \1252 , \1250 , \1251 );
mnot \mul_18_12_g22442/U$4 ( \1253 , \1250 );
mand \mul_18_12_g22442/U$3 ( \1254 , \1253 , \1198 );
mnor \mul_18_12_g22442/U$1 ( \1255 , \1252 , \1254 );
mand \mul_18_12_g22396/U$2 ( \1256 , \1245 , \1255 );
mnot \mul_18_12_g22396/U$4 ( \1257 , \1245 );
mnot \mul_18_12_g22422/U$1 ( \1258 , \1255 );
mand \mul_18_12_g22396/U$3 ( \1259 , \1257 , \1258 );
mnor \mul_18_12_g22396/U$1 ( \1260 , \1256 , \1259 );
mxnor \g36623/U$1 ( \1261 , \1177 , \1181 );
mxor \mul_18_12_g22917/U$1 ( \1262 , \a[3] , \d[3] );
mnot \mul_18_12_g22661/U$3 ( \1263 , \1262 );
mnot \mul_18_12_g22661/U$4 ( \1264 , \962 );
mor \mul_18_12_g22661/U$2 ( \1265 , \1263 , \1264 );
mnand \mul_18_12_g22730/U$1 ( \1266 , \965 , \1219 );
mnand \mul_18_12_g22661/U$1 ( \1267 , \1265 , \1266 );
mxor \mul_18_12_g37177/U$1 ( \1268 , \a[5] , \d[1] );
mnot \mul_18_12_g22688/U$3 ( \1269 , \1268 );
mnot \mul_18_12_g22688/U$4 ( \1270 , \1065 );
mor \mul_18_12_g22688/U$2 ( \1271 , \1269 , \1270 );
mnand \mul_18_12_g22734/U$1 ( \1272 , \1173 , \d[0] );
mnand \mul_18_12_g22688/U$1 ( \1273 , \1271 , \1272 );
mnot \mul_18_12_g22587/U$2 ( \1274 , \1273 );
mnand \mul_18_12_g22783/U$1 ( \1275 , \998 , \a[0] );
mnand \mul_18_12_g22587/U$1 ( \1276 , \1274 , \1275 );
mand \mul_18_12_g22497/U$2 ( \1277 , \1267 , \1276 );
mnot \mul_18_12_g22586/U$2 ( \1278 , \1273 );
mnor \mul_18_12_g22586/U$1 ( \1279 , \1278 , \1275 );
mnor \mul_18_12_g22497/U$1 ( \1280 , \1277 , \1279 );
mxor \mul_18_12_g22388/U$4 ( \1281 , \1261 , \1280 );
mxor \mul_18_12_g23065/U$1 ( \1282 , \1237 , \1230 );
mxnor \mul_18_12_g23065/U$1_r1 ( \1283 , \1282 , \1224 );
mand \mul_18_12_g22388/U$3 ( \1284 , \1281 , \1283 );
mand \mul_18_12_g22388/U$5 ( \1285 , \1261 , \1280 );
mor \mul_18_12_g22388/U$2 ( \1286 , \1284 , \1285 );
mnand \mul_18_12_g22337/U$1 ( \1287 , \1260 , \1286 );
mnot \mul_18_12_g22315/U$2 ( \1288 , \1287 );
mnot \mul_18_12_g22367/U$3 ( \1289 , \1217 );
mnot \mul_18_12_g22367/U$4 ( \1290 , \1258 );
mor \mul_18_12_g22367/U$2 ( \1291 , \1289 , \1290 );
mnot \g37119/U$3 ( \1292 , \1255 );
mnot \g37119/U$4 ( \1293 , \1216 );
mor \g37119/U$2 ( \1294 , \1292 , \1293 );
mnand \g37119/U$1 ( \1295 , \1294 , \1240 );
mnand \mul_18_12_g22367/U$1 ( \1296 , \1291 , \1295 );
mnot \mul_18_12_g22395/U$3 ( \1297 , \1202 );
mnot \mul_18_12_g22395/U$4 ( \1298 , \1170 );
mor \mul_18_12_g22395/U$2 ( \1299 , \1297 , \1298 );
mor \mul_18_12_g22395/U$5 ( \1300 , \1202 , \1170 );
mnand \mul_18_12_g22395/U$1 ( \1301 , \1299 , \1300 );
mnot \mul_18_12_g22373/U$1 ( \1302 , \1301 );
mnot \mul_18_12_g22352/U$3 ( \1303 , \1302 );
mnot \mul_18_12_g22352/U$4 ( \1304 , \1207 );
mor \mul_18_12_g22352/U$2 ( \1305 , \1303 , \1304 );
mnand \mul_18_12_g22354/U$1 ( \1306 , \1206 , \1301 );
mnand \mul_18_12_g22352/U$1 ( \1307 , \1305 , \1306 );
mnor \mul_18_12_g22325/U$1 ( \1308 , \1296 , \1307 );
mnor \mul_18_12_g22315/U$1 ( \1309 , \1288 , \1308 );
mand \mul_18_12_g23021/U$1 ( \1310 , \1161 , \1214 , \1309 );
mnot \mul_18_12_g22640/U$3 ( \1311 , \937 );
mbuf \mul_18_12_g22721/U$1 ( \1312 , \933 );
mnot \mul_18_12_g22640/U$4 ( \1313 , \1312 );
mor \mul_18_12_g22640/U$2 ( \1314 , \1311 , \1313 );
mxor \mul_18_12_g22885/U$1 ( \1315 , \a[8] , \d[5] );
mnand \mul_18_12_g22712/U$1 ( \1316 , \936 , \1315 );
mnand \mul_18_12_g22640/U$1 ( \1317 , \1314 , \1316 );
mand \mul_18_12_g22527/U$2 ( \1318 , \956 , \968 );
mxor \mul_18_12_g22412/U$1 ( \1319 , \1317 , \1318 );
mnot \mul_18_12_g22522/U$3 ( \1320 , \1096 );
mnot \mul_18_12_g22522/U$4 ( \1321 , \1117 );
mor \mul_18_12_g22522/U$2 ( \1322 , \1320 , \1321 );
mnand \mul_18_12_g22522/U$1 ( \1323 , \1322 , \1103 );
mnand \mul_18_12_g22529/U$1 ( \1324 , \1095 , \1118 );
mnand \mul_18_12_g22498/U$1 ( \1325 , \1323 , \1324 );
mxor \mul_18_12_g22412/U$1_r1 ( \1326 , \1319 , \1325 );
mbuf \mul_18_12_g22444/U$1 ( \1327 , \1081 );
mnot \mul_18_12_g22384/U$3 ( \1328 , \1327 );
mnot \mul_18_12_g22384/U$4 ( \1329 , \1124 );
mor \mul_18_12_g22384/U$2 ( \1330 , \1328 , \1329 );
mor \mul_18_12_g22406/U$2 ( \1331 , \1124 , \1327 );
mnand \mul_18_12_g22406/U$1 ( \1332 , \1331 , \1088 );
mnand \mul_18_12_g22384/U$1 ( \1333 , \1330 , \1332 );
mxor \mul_18_12_g22310/U$1 ( \1334 , \1326 , \1333 );
mxor \mul_18_12_g36683/U$1 ( \1335 , \d[12] , \d[11] );
mand \mul_18_12_g23027/U$1 ( \1336 , \1335 , \a[0] );
mnot \mul_18_12_g22624/U$3 ( \1337 , \1101 );
mnot \mul_18_12_g22624/U$4 ( \1338 , \1038 );
mor \mul_18_12_g22624/U$2 ( \1339 , \1337 , \1338 );
mxor \mul_18_12_g22899/U$1 ( \1340 , \a[6] , \d[7] );
mnand \mul_18_12_g22744/U$1 ( \1341 , \998 , \1340 );
mnand \mul_18_12_g22624/U$1 ( \1342 , \1339 , \1341 );
mxor \mul_18_12_g22454/U$1 ( \1343 , \1336 , \1342 );
mnot \mul_18_12_g22655/U$3 ( \1344 , \966 );
mnot \mul_18_12_g22655/U$4 ( \1345 , \980 );
mor \mul_18_12_g22655/U$2 ( \1346 , \1344 , \1345 );
mxor \mul_18_12_g22856/U$1 ( \1347 , \a[10] , \d[3] );
mnand \mul_18_12_g22743/U$1 ( \1348 , \965 , \1347 );
mnand \mul_18_12_g22655/U$1 ( \1349 , \1346 , \1348 );
mxor \mul_18_12_g22454/U$1_r1 ( \1350 , \1343 , \1349 );
mnot \g37124/U$3 ( \1351 , \1109 );
mnot \g37124/U$4 ( \1352 , \1115 );
mor \g37124/U$2 ( \1353 , \1351 , \1352 );
mxnor \mul_18_12_g23033/U$1 ( \1354 , \a[4] , \d[9] );
mnot \mul_18_12_g22672/U$2 ( \1355 , \1354 );
mnand \mul_18_12_g22672/U$1 ( \1356 , \1355 , \1029 );
mnand \g37124/U$1 ( \1357 , \1353 , \1356 );
mnot \mul_18_12_g22704/U$3 ( \1358 , \1065 );
mnot \mul_18_12_g22704/U$4 ( \1359 , \1093 );
mor \mul_18_12_g22704/U$2 ( \1360 , \1358 , \1359 );
mxor \g36628/U$1 ( \1361 , \d[1] , \a[12] );
mnand \mul_18_12_g22780/U$1 ( \1362 , \1361 , \d[0] );
mnand \mul_18_12_g22704/U$1 ( \1363 , \1360 , \1362 );
mxor \mul_18_12_g22510/U$1 ( \1364 , \1357 , \1363 );
mnot \mul_18_12_g22619/U$3 ( \1365 , \948 );
mnor \mul_18_12_g22812/U$1 ( \1366 , \947 , \942 );
mnot \mul_18_12_g22619/U$4 ( \1367 , \1366 );
mor \mul_18_12_g22619/U$2 ( \1368 , \1365 , \1367 );
mxor \mul_18_12_g22940/U$1 ( \1369 , \a[2] , \d[11] );
mnand \mul_18_12_g22748/U$1 ( \1370 , \947 , \1369 );
mnand \mul_18_12_g22619/U$1 ( \1371 , \1368 , \1370 );
mxor \mul_18_12_g36761/U$1 ( \1372 , \1364 , \1371 );
mxor \mul_18_12_g22350/U$1 ( \1373 , \1350 , \1372 );
mnot \mul_18_12_g22550/U$2 ( \1374 , \939 );
mnand \mul_18_12_g22550/U$1 ( \1375 , \1374 , \951 );
mnot \mul_18_12_g22472/U$3 ( \1376 , \1375 );
mnot \mul_18_12_g22472/U$4 ( \1377 , \969 );
mor \mul_18_12_g22472/U$2 ( \1378 , \1376 , \1377 );
mnand \mul_18_12_g22557/U$1 ( \1379 , \939 , \950 );
mnand \mul_18_12_g22472/U$1 ( \1380 , \1378 , \1379 );
mxor \mul_18_12_g22350/U$1_r1 ( \1381 , \1373 , \1380 );
mxor \mul_18_12_g22310/U$1_r1 ( \1382 , \1334 , \1381 );
mnor \mul_18_12_g22360/U$1 ( \1383 , \1050 , \970 );
mor \mul_18_12_g22332/U$2 ( \1384 , \1125 , \1383 );
mnand \mul_18_12_g22365/U$1 ( \1385 , \1050 , \970 );
mnand \mul_18_12_g22332/U$1 ( \1386 , \1384 , \1385 );
mnor \mul_18_12_g22292/U$1 ( \1387 , \1382 , \1386 );
mnot \mul_18_12_g22291/U$1 ( \1388 , \1387 );
mxor \mul_18_12_g22388/U$1 ( \1389 , \1261 , \1280 );
mxor \mul_18_12_g22388/U$1_r1 ( \1390 , \1389 , \1283 );
mxor \mul_18_12_g22507/U$1 ( \1391 , \1275 , \1273 );
mxnor \mul_18_12_g22507/U$1_r1 ( \1392 , \1391 , \1267 );
mor \mul_18_12_g22821/U$2 ( \1393 , \a[0] , \d[4] );
mnand \mul_18_12_g22821/U$1 ( \1394 , \1393 , \d[3] );
mnand \mul_18_12_g22961/U$1 ( \1395 , \a[0] , \d[4] );
mnand \mul_18_12_g22795/U$1 ( \1396 , \1394 , \1395 , \d[5] );
mnot \mul_18_12_g23071/U$2 ( \1397 , \1396 );
mxor \mul_18_12_g22902/U$1 ( \1398 , \a[4] , \d[1] );
mnot \mul_18_12_g22687/U$3 ( \1399 , \1398 );
mnot \mul_18_12_g22687/U$4 ( \1400 , \1012 );
mor \mul_18_12_g22687/U$2 ( \1401 , \1399 , \1400 );
mnand \mul_18_12_g22728/U$1 ( \1402 , \1268 , \d[0] );
mnand \mul_18_12_g22687/U$1 ( \1403 , \1401 , \1402 );
mnand \mul_18_12_g23071/U$1 ( \1404 , \1397 , \1403 );
mxor \mul_18_12_g22931/U$1 ( \1405 , \a[1] , \d[5] );
mnot \mul_18_12_g22647/U$3 ( \1406 , \1405 );
mnot \mul_18_12_g22647/U$4 ( \1407 , \1186 );
mor \mul_18_12_g22647/U$2 ( \1408 , \1406 , \1407 );
mnand \mul_18_12_g22765/U$1 ( \1409 , \936 , \1225 );
mnand \mul_18_12_g22647/U$1 ( \1410 , \1408 , \1409 );
mnot \mul_18_12_g22646/U$1 ( \1411 , \1410 );
mnand \mul_18_12_g22515/U$1 ( \1412 , \1404 , \1411 );
mand \mul_18_12_g22435/U$2 ( \1413 , \1392 , \1412 );
mnot \mul_18_12_g22543/U$1 ( \1414 , \1404 );
mand \mul_18_12_g23022/U$1 ( \1415 , \1414 , \1410 );
mnor \mul_18_12_g22435/U$1 ( \1416 , \1413 , \1415 );
mnand \mul_18_12_g22364/U$1 ( \1417 , \1390 , \1416 );
mnot \mul_18_12_g22279/U$3 ( \1418 , \1417 );
mnot \mul_18_12_g22597/U$3 ( \1419 , \1405 );
mnot \mul_18_12_g22597/U$4 ( \1420 , \932 );
mor \mul_18_12_g22597/U$2 ( \1421 , \1419 , \1420 );
mxor \mul_18_12_g22945/U$1 ( \1422 , \a[0] , \d[5] );
mnand \mul_18_12_g22741/U$1 ( \1423 , \930 , \1422 );
mor \mul_18_12_g22597/U$5 ( \1424 , \932 , \1423 );
mnand \mul_18_12_g22597/U$1 ( \1425 , \1421 , \1424 );
mxor \mul_18_12_g37178/U$1 ( \1426 , \a[2] , \d[3] );
mnot \mul_18_12_g22665/U$3 ( \1427 , \1426 );
mnot \mul_18_12_g22665/U$4 ( \1428 , \980 );
mor \mul_18_12_g22665/U$2 ( \1429 , \1427 , \1428 );
mnand \mul_18_12_g22753/U$1 ( \1430 , \965 , \1262 );
mnand \mul_18_12_g22665/U$1 ( \1431 , \1429 , \1430 );
mxor \mul_18_12_g22426/U$4 ( \1432 , \1425 , \1431 );
mnot \mul_18_12_g22577/U$3 ( \1433 , \1396 );
mnot \mul_18_12_g22577/U$4 ( \1434 , \1403 );
mor \mul_18_12_g22577/U$2 ( \1435 , \1433 , \1434 );
mor \mul_18_12_g22577/U$5 ( \1436 , \1403 , \1396 );
mnand \mul_18_12_g22577/U$1 ( \1437 , \1435 , \1436 );
mand \mul_18_12_g22426/U$3 ( \1438 , \1432 , \1437 );
mand \mul_18_12_g22426/U$5 ( \1439 , \1425 , \1431 );
mor \mul_18_12_g22426/U$2 ( \1440 , \1438 , \1439 );
mxor \g36621/U$1 ( \1441 , \1414 , \1411 );
mxnor \g36621/U$1_r1 ( \1442 , \1441 , \1392 );
mxor \mul_18_12_g22308/U$4 ( \1443 , \1440 , \1442 );
mxor \mul_18_12_g22426/U$1 ( \1444 , \1425 , \1431 );
mxor \mul_18_12_g22426/U$1_r1 ( \1445 , \1444 , \1437 );
mxor \mul_18_12_g22929/U$1 ( \1446 , \a[1] , \d[3] );
mnand \mul_18_12_g22767/U$1 ( \1447 , \961 , \1446 );
mor \mul_18_12_g22600/U$2 ( \1448 , \1447 , \965 );
mnand \mul_18_12_g22747/U$1 ( \1449 , \959 , \1426 );
mnand \mul_18_12_g22600/U$1 ( \1450 , \1448 , \1449 );
mnot \g37122/U$3 ( \1451 , \1450 );
mxor \g36636/U$1 ( \1452 , \d[1] , \a[3] );
mnot \mul_18_12_g22690/U$3 ( \1453 , \1452 );
mnot \mul_18_12_g22690/U$4 ( \1454 , \1012 );
mor \mul_18_12_g22690/U$2 ( \1455 , \1453 , \1454 );
mnand \mul_18_12_g22758/U$1 ( \1456 , \1398 , \d[0] );
mnand \mul_18_12_g22690/U$1 ( \1457 , \1455 , \1456 );
mnot \mul_18_12_g22589/U$2 ( \1458 , \1457 );
mnand \mul_18_12_g22786/U$1 ( \1459 , \932 , \a[0] );
mnand \mul_18_12_g22589/U$1 ( \1460 , \1458 , \1459 );
mnot \g37122/U$4 ( \1461 , \1460 );
mor \g37122/U$2 ( \1462 , \1451 , \1461 );
mnot \mul_18_12_g23070/U$2 ( \1463 , \1459 );
mnand \mul_18_12_g23070/U$1 ( \1464 , \1463 , \1457 );
mnand \g37122/U$1 ( \1465 , \1462 , \1464 );
mnor \mul_18_12_g22401/U$1 ( \1466 , \1445 , \1465 );
mxor \g36637/U$1 ( \1467 , \d[1] , \a[2] );
mand \g37129/U$2 ( \1468 , \1065 , \1467 );
mand \g37129/U$3 ( \1469 , \1452 , \d[0] );
mnor \g37129/U$1 ( \1470 , \1468 , \1469 );
mor \mul_18_12_g22822/U$2 ( \1471 , \a[0] , \d[2] );
mnand \mul_18_12_g22822/U$1 ( \1472 , \1471 , \d[1] );
mnand \mul_18_12_g22958/U$1 ( \1473 , \a[0] , \d[2] );
mnand \mul_18_12_g22793/U$1 ( \1474 , \1472 , \1473 , \d[3] );
mnot \mul_18_12_g22792/U$1 ( \1475 , \1474 );
mand \mul_18_12_g22578/U$2 ( \1476 , \1470 , \1475 );
mnot \mul_18_12_g22578/U$4 ( \1477 , \1470 );
mand \mul_18_12_g22578/U$3 ( \1478 , \1477 , \1474 );
mnor \mul_18_12_g22578/U$1 ( \1479 , \1476 , \1478 );
mnot \mul_18_12_g22602/U$3 ( \1480 , \965 );
mxor \mul_18_12_g22949/U$1 ( \1481 , \a[0] , \d[3] );
mnand \mul_18_12_g22755/U$1 ( \1482 , \961 , \1481 );
mnot \mul_18_12_g22602/U$4 ( \1483 , \1482 );
mand \mul_18_12_g22602/U$2 ( \1484 , \1480 , \1483 );
mand \mul_18_12_g22602/U$5 ( \1485 , \965 , \1446 );
mnor \mul_18_12_g22602/U$1 ( \1486 , \1484 , \1485 );
mor \mul_18_12_g23056/U$1 ( \1487 , \1479 , \1486 );
mnand \mul_18_12_g22519/U$1 ( \1488 , \1479 , \1486 );
mxor \g36638/U$1 ( \1489 , \d[1] , \a[1] );
mnot \mul_18_12_g22693/U$3 ( \1490 , \1489 );
mnot \mul_18_12_g22693/U$4 ( \1491 , \1012 );
mor \mul_18_12_g22693/U$2 ( \1492 , \1490 , \1491 );
mnand \mul_18_12_g22708/U$1 ( \1493 , \1467 , \d[0] );
mnand \mul_18_12_g22693/U$1 ( \1494 , \1492 , \1493 );
mand \mul_18_12_g23028/U$1 ( \1495 , \959 , \a[0] );
mnor \mul_18_12_g22590/U$1 ( \1496 , \1494 , \1495 );
mxor \mul_18_12_g22950/U$1 ( \1497 , \a[0] , \d[1] );
mnot \mul_18_12_g22697/U$3 ( \1498 , \1497 );
mnot \mul_18_12_g22697/U$4 ( \1499 , \1012 );
mor \mul_18_12_g22697/U$2 ( \1500 , \1498 , \1499 );
mnand \mul_18_12_g22757/U$1 ( \1501 , \1489 , \d[0] );
mnand \mul_18_12_g22697/U$1 ( \1502 , \1500 , \1501 );
mand \mul_18_12_g22815/U$1 ( \1503 , \684 , \d[1] );
mnand \mul_18_12_g22585/U$1 ( \1504 , \1502 , \1503 );
mor \mul_18_12_g22496/U$2 ( \1505 , \1496 , \1504 );
mnand \mul_18_12_g22591/U$1 ( \1506 , \1494 , \1495 );
mnand \mul_18_12_g22496/U$1 ( \1507 , \1505 , \1506 );
mnand \mul_18_12_g22449/U$1 ( \1508 , \1488 , \1507 );
mnand \mul_18_12_g22434/U$1 ( \1509 , \1487 , \1508 );
mxor \g36906/U$1 ( \1510 , \1459 , \1450 );
mxor \g36906/U$1_r1 ( \1511 , \1510 , \1457 );
mnot \mul_18_12_g23067/U$2 ( \1512 , \1470 );
mnand \mul_18_12_g23067/U$1 ( \1513 , \1512 , \1475 );
mnand \mul_18_12_g22448/U$1 ( \1514 , \1511 , \1513 );
mand \mul_18_12_g22381/U$2 ( \1515 , \1509 , \1514 );
mnor \mul_18_12_g22447/U$1 ( \1516 , \1511 , \1513 );
mnor \mul_18_12_g22381/U$1 ( \1517 , \1515 , \1516 );
mor \mul_18_12_g22340/U$2 ( \1518 , \1466 , \1517 );
mnand \mul_18_12_g22400/U$1 ( \1519 , \1445 , \1465 );
mnand \mul_18_12_g22340/U$1 ( \1520 , \1518 , \1519 );
mand \mul_18_12_g22308/U$3 ( \1521 , \1443 , \1520 );
mand \mul_18_12_g22308/U$5 ( \1522 , \1440 , \1442 );
mor \mul_18_12_g22308/U$2 ( \1523 , \1521 , \1522 );
mnot \mul_18_12_g22279/U$4 ( \1524 , \1523 );
mor \mul_18_12_g22279/U$2 ( \1525 , \1418 , \1524 );
mor \g37070/U$1 ( \1526 , \1390 , \1416 );
mnand \mul_18_12_g22279/U$1 ( \1527 , \1525 , \1526 );
mbuf \mul_18_12_g22268/U$1 ( \1528 , \1527 );
mnand \mul_18_12_g22252/U$1 ( \1529 , \1310 , \1388 , \1528 );
mnor \mul_18_12_g22289/U$1 ( \1530 , \1160 , \1126 );
mnand \g36612/U$1 ( \1531 , \1388 , \1530 );
mnot \mul_18_12_g22358/U$1 ( \1532 , \1260 );
mnot \mul_18_12_g22387/U$1 ( \1533 , \1286 );
mnand \mul_18_12_g22339/U$1 ( \1534 , \1532 , \1533 );
mor \mul_18_12_g22305/U$2 ( \1535 , \1308 , \1534 );
mnand \mul_18_12_g22324/U$1 ( \1536 , \1307 , \1296 );
mnand \mul_18_12_g22305/U$1 ( \1537 , \1535 , \1536 );
mnor \mul_18_12_g22318/U$1 ( \1538 , \1163 , \1213 );
mnor \mul_18_12_g22293/U$1 ( \1539 , \1537 , \1538 );
mnot \mul_18_12_g22267/U$2 ( \1540 , \1539 );
mbuf \mul_18_12_g22286/U$1 ( \1541 , \1161 );
mnand \mul_18_12_g22267/U$1 ( \1542 , \1540 , \1541 , \1214 , \1388 );
mnand \mul_18_12_g22297/U$1 ( \1543 , \1382 , \1386 );
mnand \mul_18_12_g22241/U$1 ( \1544 , \1529 , \1531 , \1542 , \1543 );
mnot \mul_18_12_g22700/U$3 ( \1545 , \1361 );
mnot \mul_18_12_g22700/U$4 ( \1546 , \1065 );
mor \mul_18_12_g22700/U$2 ( \1547 , \1545 , \1546 );
mxor \mul_18_12_g22843/U$1 ( \1548 , \a[13] , \d[1] );
mnand \mul_18_12_g22778/U$1 ( \1549 , \1548 , \d[0] );
mnand \mul_18_12_g22700/U$1 ( \1550 , \1547 , \1549 );
mnot \mul_18_12_g22560/U$3 ( \1551 , \1550 );
mor \mul_18_12_g22817/U$2 ( \1552 , \a[0] , \d[12] );
mnand \mul_18_12_g22817/U$1 ( \1553 , \1552 , \d[11] );
mnand \mul_18_12_g22957/U$1 ( \1554 , \a[0] , \d[12] );
mnand \mul_18_12_g22805/U$1 ( \1555 , \1553 , \1554 , \d[13] );
mnot \mul_18_12_g22560/U$4 ( \1556 , \1555 );
mand \mul_18_12_g22560/U$2 ( \1557 , \1551 , \1556 );
mand \mul_18_12_g22560/U$5 ( \1558 , \1550 , \1555 );
mnor \mul_18_12_g22560/U$1 ( \1559 , \1557 , \1558 );
mxor \mul_18_12_g22454/U$4 ( \1560 , \1336 , \1342 );
mand \mul_18_12_g22454/U$3 ( \1561 , \1560 , \1349 );
mand \mul_18_12_g22454/U$5 ( \1562 , \1336 , \1342 );
mor \mul_18_12_g22454/U$2 ( \1563 , \1561 , \1562 );
mxor \mul_18_12_g36786/U$1 ( \1564 , \1559 , \1563 );
mor \mul_18_12_g23057/U$1 ( \1565 , \1357 , \1363 );
mand \mul_18_12_g22452/U$2 ( \1566 , \1565 , \1371 );
mand \mul_18_12_g22510/U$2 ( \1567 , \1357 , \1363 );
mnor \mul_18_12_g22452/U$1 ( \1568 , \1566 , \1567 );
mnot \mul_18_12_g22443/U$1 ( \1569 , \1568 );
mxor \mul_18_12_g36786/U$1_r1 ( \1570 , \1564 , \1569 );
mnot \mul_18_12_g22329/U$3 ( \1571 , \1570 );
mxor \mul_18_12_g22350/U$4 ( \1572 , \1350 , \1372 );
mand \mul_18_12_g22350/U$3 ( \1573 , \1572 , \1380 );
mand \mul_18_12_g22350/U$5 ( \1574 , \1350 , \1372 );
mor \mul_18_12_g22350/U$2 ( \1575 , \1573 , \1574 );
mnot \mul_18_12_g22329/U$4 ( \1576 , \1575 );
mor \mul_18_12_g22329/U$2 ( \1577 , \1571 , \1576 );
mor \mul_18_12_g22329/U$5 ( \1578 , \1575 , \1570 );
mnand \mul_18_12_g22329/U$1 ( \1579 , \1577 , \1578 );
mxor \mul_18_12_g22913/U$1 ( \1580 , \a[0] , \d[13] );
mnot \mul_18_12_g22609/U$3 ( \1581 , \1580 );
mxnor \mul_18_12_g23031/U$1 ( \1582 , \d[13] , \d[12] );
mnor \mul_18_12_g22809/U$1 ( \1583 , \1582 , \1335 );
mnot \mul_18_12_g22609/U$4 ( \1584 , \1583 );
mor \mul_18_12_g22609/U$2 ( \1585 , \1581 , \1584 );
mxor \mul_18_12_g22942/U$1 ( \1586 , \a[1] , \d[13] );
mnand \mul_18_12_g22713/U$1 ( \1587 , \1335 , \1586 );
mnand \mul_18_12_g22609/U$1 ( \1588 , \1585 , \1587 );
mnot \mul_18_12_g22620/U$3 ( \1589 , \1369 );
mnot \mul_18_12_g22620/U$4 ( \1590 , \944 );
mor \mul_18_12_g22620/U$2 ( \1591 , \1589 , \1590 );
mxor \mul_18_12_g22939/U$1 ( \1592 , \a[3] , \d[11] );
mnand \mul_18_12_g22766/U$1 ( \1593 , \947 , \1592 );
mnand \mul_18_12_g22620/U$1 ( \1594 , \1591 , \1593 );
mxor \mul_18_12_g22484/U$1 ( \1595 , \1588 , \1594 );
mnot \mul_18_12_g22653/U$3 ( \1596 , \1315 );
mnot \mul_18_12_g22653/U$4 ( \1597 , \933 );
mor \mul_18_12_g22653/U$2 ( \1598 , \1596 , \1597 );
mxor \mul_18_12_g22884/U$1 ( \1599 , \a[9] , \d[5] );
mnand \mul_18_12_g22764/U$1 ( \1600 , \936 , \1599 );
mnand \mul_18_12_g22653/U$1 ( \1601 , \1598 , \1600 );
mxor \mul_18_12_g22484/U$1_r1 ( \1602 , \1595 , \1601 );
mnot \mul_18_12_g22483/U$1 ( \1603 , \1602 );
mnot \mul_18_12_g22428/U$3 ( \1604 , \1603 );
mnot \mul_18_12_g22570/U$3 ( \1605 , \1110 );
mnot \mul_18_12_g22570/U$4 ( \1606 , \1354 );
mand \mul_18_12_g22570/U$2 ( \1607 , \1605 , \1606 );
mxor \mul_18_12_g37176/U$1 ( \1608 , \a[5] , \d[9] );
mand \mul_18_12_g22570/U$5 ( \1609 , \1058 , \1608 );
mnor \mul_18_12_g22570/U$1 ( \1610 , \1607 , \1609 );
mnot \fopt36733/U$1 ( \1611 , \1610 );
mnot \mul_18_12_g22524/U$3 ( \1612 , \1611 );
mnot \mul_18_12_g22634/U$3 ( \1613 , \1340 );
mnot \mul_18_12_g22634/U$4 ( \1614 , \999 );
mor \mul_18_12_g22634/U$2 ( \1615 , \1613 , \1614 );
mxor \mul_18_12_g22898/U$1 ( \1616 , \a[7] , \d[7] );
mnand \mul_18_12_g22754/U$1 ( \1617 , \1003 , \1616 );
mnand \mul_18_12_g22634/U$1 ( \1618 , \1615 , \1617 );
mnot \mul_18_12_g22633/U$1 ( \1619 , \1618 );
mnot \mul_18_12_g22524/U$4 ( \1620 , \1619 );
mor \mul_18_12_g22524/U$2 ( \1621 , \1612 , \1620 );
mnand \mul_18_12_g22530/U$1 ( \1622 , \1610 , \1618 );
mnand \mul_18_12_g22524/U$1 ( \1623 , \1621 , \1622 );
mnot \mul_18_12_g22657/U$3 ( \1624 , \1347 );
mnot \mul_18_12_g22657/U$4 ( \1625 , \962 );
mor \mul_18_12_g22657/U$2 ( \1626 , \1624 , \1625 );
mxor \mul_18_12_g22857/U$1 ( \1627 , \a[11] , \d[3] );
mnand \mul_18_12_g22750/U$1 ( \1628 , \965 , \1627 );
mnand \mul_18_12_g22657/U$1 ( \1629 , \1626 , \1628 );
mxnor \mul_18_12_g23064/U$1 ( \1630 , \1623 , \1629 );
mnot \mul_18_12_g22457/U$1 ( \1631 , \1630 );
mnot \mul_18_12_g22428/U$4 ( \1632 , \1631 );
mor \mul_18_12_g22428/U$2 ( \1633 , \1604 , \1632 );
mnand \mul_18_12_g22430/U$1 ( \1634 , \1630 , \1602 );
mnand \mul_18_12_g22428/U$1 ( \1635 , \1633 , \1634 );
mxor \mul_18_12_g22412/U$4 ( \1636 , \1317 , \1318 );
mand \mul_18_12_g22412/U$3 ( \1637 , \1636 , \1325 );
mand \mul_18_12_g22412/U$5 ( \1638 , \1317 , \1318 );
mor \mul_18_12_g22412/U$2 ( \1639 , \1637 , \1638 );
mnot \mul_18_12_g22411/U$1 ( \1640 , \1639 );
mand \mul_18_12_g22375/U$2 ( \1641 , \1635 , \1640 );
mnot \mul_18_12_g22375/U$4 ( \1642 , \1635 );
mand \mul_18_12_g22375/U$3 ( \1643 , \1642 , \1639 );
mnor \mul_18_12_g22375/U$1 ( \1644 , \1641 , \1643 );
mand \mul_18_12_g22311/U$2 ( \1645 , \1579 , \1644 );
mnot \mul_18_12_g22311/U$4 ( \1646 , \1579 );
mnot \mul_18_12_g22346/U$1 ( \1647 , \1644 );
mand \mul_18_12_g22311/U$3 ( \1648 , \1646 , \1647 );
mnor \mul_18_12_g22311/U$1 ( \1649 , \1645 , \1648 );
mnot \mul_18_12_g23037/U$2 ( \1650 , \1649 );
mxor \mul_18_12_g22310/U$4 ( \1651 , \1326 , \1333 );
mand \mul_18_12_g22310/U$3 ( \1652 , \1651 , \1381 );
mand \mul_18_12_g22310/U$5 ( \1653 , \1326 , \1333 );
mor \mul_18_12_g22310/U$2 ( \1654 , \1652 , \1653 );
mnand \mul_18_12_g23037/U$1 ( \1655 , \1650 , \1654 );
mnot \mul_18_12_g22274/U$2 ( \1656 , \1654 );
mnand \mul_18_12_g22274/U$1 ( \1657 , \1656 , \1649 );
mnand \mul_18_12_g22263/U$1 ( \1658 , \1655 , \1657 );
mnot \mul_18_12_g22262/U$1 ( \1659 , \1658 );
mand \mul_18_12_g22236/U$2 ( \1660 , \1544 , \1659 );
mnot \mul_18_12_g22236/U$4 ( \1661 , \1544 );
mand \mul_18_12_g22236/U$3 ( \1662 , \1661 , \1658 );
mnor \mul_18_12_g22236/U$1 ( \1663 , \1660 , \1662 );
mnand \mul_6_11_g6543/U$1 ( \1664 , \239 , \343 );
mbuf \mul_6_11_g6531/U$1 ( \1665 , \339 );
mxnor \mul_6_11_g6915/U$1 ( \1666 , \1664 , \1665 );
mnot \g4879/U$1 ( \1667 , \1666 );
mnot \g4873/U$1 ( \1668 , \1667 );
mnand \g4750/U$1 ( \1669 , \1663 , \1668 );
mxor \g36595/U$1 ( \1670 , \c[5] , \b[6] );
mnot \mul_19_13_g22638/U$3 ( \1671 , \1670 );
mxor \mul_19_13_g22870/U$1 ( \1672 , \c[5] , \c[4] );
mnot \mul_19_13_g22722/U$2 ( \1673 , \1672 );
mxor \mul_19_13_g36674/U$1 ( \1674 , \c[4] , \c[3] );
mnor \mul_19_13_g22722/U$1 ( \1675 , \1673 , \1674 );
mnot \mul_19_13_g22638/U$4 ( \1676 , \1675 );
mor \mul_19_13_g22638/U$2 ( \1677 , \1671 , \1676 );
mbuf \mul_19_13_g22851/U$1 ( \1678 , \1674 );
mxor \g36594/U$1 ( \1679 , \c[5] , \b[7] );
mnand \mul_19_13_g22710/U$1 ( \1680 , \1678 , \1679 );
mnand \mul_19_13_g22638/U$1 ( \1681 , \1677 , \1680 );
mxor \mul_19_13_g22930/U$1 ( \1682 , \b[0] , \c[11] );
mnot \mul_19_13_g22615/U$3 ( \1683 , \1682 );
mxnor \mul_19_13_g36687/U$1 ( \1684 , \c[11] , \c[10] );
mxor \mul_19_13_g22875/U$1 ( \1685 , \c[10] , \c[9] );
mnor \mul_19_13_g22811/U$1 ( \1686 , \1684 , \1685 );
mnot \mul_19_13_g22615/U$4 ( \1687 , \1686 );
mor \mul_19_13_g22615/U$2 ( \1688 , \1683 , \1687 );
mxor \mul_19_13_g22876/U$1 ( \1689 , \c[10] , \c[9] );
mxor \mul_19_13_g22944/U$1 ( \1690 , \b[1] , \c[11] );
mnand \mul_19_13_g22711/U$1 ( \1691 , \1689 , \1690 );
mnand \mul_19_13_g22615/U$1 ( \1692 , \1688 , \1691 );
mnot \mul_19_13_g22614/U$1 ( \1693 , \1692 );
mxor \g36578/U$1 ( \1694 , \1681 , \1693 );
mor \mul_19_13_g22818/U$2 ( \1695 , \b[0] , \c[10] );
mnand \mul_19_13_g22818/U$1 ( \1696 , \1695 , \c[9] );
mnand \mul_19_13_g22956/U$1 ( \1697 , \b[0] , \c[10] );
mand \mul_19_13_g23029/U$1 ( \1698 , \1696 , \1697 , \c[11] );
mxor \mul_19_13_g22883/U$1 ( \1699 , \b[8] , \c[3] );
mnot \mul_19_13_g22662/U$3 ( \1700 , \1699 );
mxor \mul_19_13_g22855/U$1 ( \1701 , \c[3] , \c[2] );
mbuf \mul_19_13_g22854/U$1 ( \1702 , \1701 );
mxor \mul_19_13_g23018/U$1 ( \1703 , \c[2] , \c[1] );
mnot \fopt37002/U$1 ( \1704 , \1703 );
mand \mul_19_13_g22761/U$1 ( \1705 , \1702 , \1704 );
mnot \mul_19_13_g22662/U$4 ( \1706 , \1705 );
mor \mul_19_13_g22662/U$2 ( \1707 , \1700 , \1706 );
mbuf \fopt37000/U$1 ( \1708 , \1703 );
mxor \mul_19_13_g22882/U$1 ( \1709 , \b[9] , \c[3] );
mnand \mul_19_13_g22729/U$1 ( \1710 , \1708 , \1709 );
mnand \mul_19_13_g22662/U$1 ( \1711 , \1707 , \1710 );
mxor \mul_19_13_g22527/U$1 ( \1712 , \1698 , \1711 );
mxnor \g36578/U$1_r1 ( \1713 , \1694 , \1712 );
mor \mul_19_13_g22819/U$2 ( \1714 , \b[0] , \c[8] );
mnand \mul_19_13_g22819/U$1 ( \1715 , \1714 , \c[7] );
mnand \mul_19_13_g22951/U$1 ( \1716 , \b[0] , \c[8] );
mnand \mul_19_13_g22799/U$1 ( \1717 , \1715 , \1716 , \c[9] );
mnot \mul_19_13_g23072/U$2 ( \1718 , \1717 );
mxor \mul_19_13_g22895/U$1 ( \1719 , \b[6] , \c[3] );
mnot \mul_19_13_g22666/U$3 ( \1720 , \1719 );
mnot \mul_19_13_g22760/U$2 ( \1721 , \1701 );
mnor \mul_19_13_g22760/U$1 ( \1722 , \1721 , \1703 );
mnot \mul_19_13_g22666/U$4 ( \1723 , \1722 );
mor \mul_19_13_g22666/U$2 ( \1724 , \1720 , \1723 );
mnot \fopt37001/U$1 ( \1725 , \1704 );
mxor \mul_19_13_g22893/U$1 ( \1726 , \b[7] , \c[3] );
mnand \mul_19_13_g22732/U$1 ( \1727 , \1725 , \1726 );
mnand \mul_19_13_g22666/U$1 ( \1728 , \1724 , \1727 );
mnand \mul_19_13_g23072/U$1 ( \1729 , \1718 , \1728 );
mnot \mul_19_13_g22416/U$3 ( \1730 , \1729 );
mnand \mul_19_13_g36688/U$1 ( \1731 , \1685 , \b[0] );
mnot \mul_19_13_g22776/U$1 ( \1732 , \1731 );
mand \g36588/U$2 ( \1733 , \1703 , \1699 );
mnot \g36588/U$4 ( \1734 , \1703 );
mand \g3/U$1 ( \1735 , \1701 , \1726 );
mand \g36588/U$3 ( \1736 , \1734 , \1735 );
mor \g36588/U$1 ( \1737 , \1733 , \1736 );
mxor \mul_19_13_g22475/U$1 ( \1738 , \1732 , \1737 );
mxor \g36601/U$1 ( \1739 , \c[7] , \b[3] );
mnot \mul_19_13_g22626/U$3 ( \1740 , \1739 );
mxnor \mul_19_13_g23032/U$1 ( \1741 , \c[7] , \c[6] );
mxor \mul_19_13_g36676/U$1 ( \1742 , \c[6] , \c[5] );
mnor \mul_19_13_g22707/U$1 ( \1743 , \1741 , \1742 );
mnot \mul_19_13_g22626/U$4 ( \1744 , \1743 );
mor \mul_19_13_g22626/U$2 ( \1745 , \1740 , \1744 );
mnot \mul_19_13_g22868/U$1 ( \1746 , \1742 );
mnot \mul_19_13_g22864/U$1 ( \1747 , \1746 );
mxor \g36596/U$1 ( \1748 , \c[7] , \b[4] );
mnand \mul_19_13_g22705/U$1 ( \1749 , \1747 , \1748 );
mnand \mul_19_13_g22626/U$1 ( \1750 , \1745 , \1749 );
mxnor \mul_19_13_g22475/U$1_r1 ( \1751 , \1738 , \1750 );
mnot \mul_19_13_g22416/U$4 ( \1752 , \1751 );
mor \mul_19_13_g22416/U$2 ( \1753 , \1730 , \1752 );
mnot \mul_19_13_g23019/U$2 ( \1754 , \c[0] );
mnand \mul_19_13_g23019/U$1 ( \1755 , \1754 , \c[1] );
mnot \mul_19_13_g22998/U$1 ( \1756 , \1755 );
mxor \g36590/U$1 ( \1757 , \c[1] , \b[8] );
mand \g37112/U$2 ( \1758 , \1756 , \1757 );
mxor \g36591/U$1 ( \1759 , \c[1] , \b[9] );
mand \g37112/U$3 ( \1760 , \1759 , \c[0] );
mnor \g37112/U$1 ( \1761 , \1758 , \1760 );
mnot \mul_19_13_g22698/U$1 ( \1762 , \1761 );
mnot \mul_19_13_g22499/U$3 ( \1763 , \1762 );
mxor \g36603/U$1 ( \1764 , \c[9] , \b[0] );
mnot \mul_19_13_g22573/U$3 ( \1765 , \1764 );
mnot \mul_19_13_g23011/U$2 ( \1766 , \c[7] );
mnand \mul_19_13_g23011/U$1 ( \1767 , \1766 , \c[8] );
mor \mul_19_13_g37019/U$1 ( \1768 , \c[9] , \c[8] );
mnand \mul_19_13_g37171/U$1 ( \1769 , \c[9] , \c[7] );
mand \mul_19_13_g22678/U$1 ( \1770 , \1767 , \1768 , \1769 );
mnot \mul_19_13_g22573/U$4 ( \1771 , \1770 );
mor \mul_19_13_g22573/U$2 ( \1772 , \1765 , \1771 );
mxor \mul_19_13_g22823/U$1 ( \1773 , \c[8] , \c[7] );
mxor \g36604/U$1 ( \1774 , \c[9] , \b[1] );
mnand \mul_19_13_g22670/U$1 ( \1775 , \1773 , \1774 );
mnand \mul_19_13_g22573/U$1 ( \1776 , \1772 , \1775 );
mnot \mul_19_13_g22499/U$4 ( \1777 , \1776 );
mor \mul_19_13_g22499/U$2 ( \1778 , \1763 , \1777 );
mor \mul_19_13_g22520/U$2 ( \1779 , \1776 , \1762 );
mxor \g36600/U$1 ( \1780 , \c[7] , \b[2] );
mnot \mul_19_13_g22622/U$3 ( \1781 , \1780 );
mnor \mul_19_13_g22706/U$1 ( \1782 , \1741 , \1742 );
mnot \mul_19_13_g22622/U$4 ( \1783 , \1782 );
mor \mul_19_13_g22622/U$2 ( \1784 , \1781 , \1783 );
mnot \mul_19_13_g23074/U$2 ( \1785 , \1746 );
mnand \mul_19_13_g23074/U$1 ( \1786 , \1785 , \1739 );
mnand \mul_19_13_g22622/U$1 ( \1787 , \1784 , \1786 );
mnand \mul_19_13_g22520/U$1 ( \1788 , \1779 , \1787 );
mnand \mul_19_13_g22499/U$1 ( \1789 , \1778 , \1788 );
mnand \mul_19_13_g22416/U$1 ( \1790 , \1753 , \1789 );
mnot \mul_19_13_g23055/U$2 ( \1791 , \1729 );
mnot \mul_19_13_g22466/U$1 ( \1792 , \1751 );
mnand \mul_19_13_g23055/U$1 ( \1793 , \1791 , \1792 );
mnand \mul_19_13_g22408/U$1 ( \1794 , \1790 , \1793 );
mxor \mul_19_13_g23046/U$1 ( \1795 , \1713 , \1794 );
mxor \mul_19_13_g22935/U$1 ( \1796 , \b[2] , \c[9] );
mnot \mul_19_13_g22571/U$3 ( \1797 , \1796 );
mnot \mul_19_13_g22824/U$3 ( \1798 , \c[7] );
mnot \mul_19_13_g23015/U$1 ( \1799 , \c[8] );
mnot \mul_19_13_g22824/U$4 ( \1800 , \1799 );
mor \mul_19_13_g22824/U$2 ( \1801 , \1798 , \1800 );
mnand \mul_19_13_g22824/U$1 ( \1802 , \1801 , \1767 );
mnot \mul_19_13_g22571/U$4 ( \1803 , \1802 );
mor \mul_19_13_g22571/U$2 ( \1804 , \1797 , \1803 );
mnand \mul_19_13_g22582/U$1 ( \1805 , \1770 , \1774 );
mnand \mul_19_13_g22571/U$1 ( \1806 , \1804 , \1805 );
mnot \mul_19_13_g22695/U$3 ( \1807 , \1759 );
mnot \mul_19_13_g22695/U$4 ( \1808 , \1756 );
mor \mul_19_13_g22695/U$2 ( \1809 , \1807 , \1808 );
mxor \mul_19_13_g22845/U$1 ( \1810 , \b[10] , \c[1] );
mnand \mul_19_13_g22749/U$1 ( \1811 , \1810 , \c[0] );
mnand \mul_19_13_g22695/U$1 ( \1812 , \1809 , \1811 );
mor \mul_19_13_g22470/U$2 ( \1813 , \1806 , \1812 );
mxor \mul_19_13_g22910/U$1 ( \1814 , \b[5] , \c[5] );
mnot \mul_19_13_g22652/U$3 ( \1815 , \1814 );
mnot \mul_19_13_g22652/U$4 ( \1816 , \1675 );
mor \mul_19_13_g22652/U$2 ( \1817 , \1815 , \1816 );
mnand \mul_19_13_g22763/U$1 ( \1818 , \1678 , \1670 );
mnand \mul_19_13_g22652/U$1 ( \1819 , \1817 , \1818 );
mnand \mul_19_13_g22470/U$1 ( \1820 , \1813 , \1819 );
mnand \mul_19_13_g22532/U$1 ( \1821 , \1806 , \1812 );
mnand \mul_19_13_g22451/U$1 ( \1822 , \1820 , \1821 );
mnot \g37162/U$2 ( \1823 , \1737 );
mnand \g37162/U$1 ( \1824 , \1823 , \1731 );
mnot \g37161/U$3 ( \1825 , \1824 );
mnot \g37161/U$4 ( \1826 , \1750 );
mor \g37161/U$2 ( \1827 , \1825 , \1826 );
mnand \mul_19_13_g22553/U$1 ( \1828 , \1737 , \1732 );
mnand \g37161/U$1 ( \1829 , \1827 , \1828 );
mxor \g37114/U$1 ( \1830 , \1822 , \1829 );
mnot \mul_19_13_g22630/U$3 ( \1831 , \1748 );
mnot \mul_19_13_g22630/U$4 ( \1832 , \1782 );
mor \mul_19_13_g22630/U$2 ( \1833 , \1831 , \1832 );
mxor \mul_19_13_g22911/U$1 ( \1834 , \b[5] , \c[7] );
mnand \mul_19_13_g22745/U$1 ( \1835 , \1747 , \1834 );
mnand \mul_19_13_g22630/U$1 ( \1836 , \1833 , \1835 );
mnot \mul_19_13_g22684/U$3 ( \1837 , \1810 );
mnot \mul_19_13_g22684/U$4 ( \1838 , \1756 );
mor \mul_19_13_g22684/U$2 ( \1839 , \1837 , \1838 );
mxor \mul_19_13_g22844/U$1 ( \1840 , \b[11] , \c[1] );
mnand \mul_19_13_g22738/U$1 ( \1841 , \1840 , \c[0] );
mnand \mul_19_13_g22684/U$1 ( \1842 , \1839 , \1841 );
mnot \mul_19_13_g22683/U$1 ( \1843 , \1842 );
mand \g37282/U$2 ( \1844 , \1836 , \1843 );
mnot \g37282/U$4 ( \1845 , \1836 );
mand \g37282/U$3 ( \1846 , \1845 , \1842 );
mor \g37282/U$1 ( \1847 , \1844 , \1846 );
mnot \mul_19_13_g22679/U$2 ( \1848 , \1767 );
mor \g37018/U$2 ( \1849 , \c[9] , \c[8] );
mnand \g37018/U$1 ( \1850 , \1849 , \1769 );
mnor \mul_19_13_g22679/U$1 ( \1851 , \1848 , \1850 );
mnot \mul_19_13_g22677/U$1 ( \1852 , \1851 );
mnot \mul_19_13_g22564/U$3 ( \1853 , \1852 );
mnot \mul_19_13_g22934/U$1 ( \1854 , \1796 );
mnot \mul_19_13_g22564/U$4 ( \1855 , \1854 );
mand \mul_19_13_g22564/U$2 ( \1856 , \1853 , \1855 );
mxor \mul_19_13_g22936/U$1 ( \1857 , \b[3] , \c[9] );
mand \mul_19_13_g22564/U$5 ( \1858 , \1802 , \1857 );
mnor \mul_19_13_g22564/U$1 ( \1859 , \1856 , \1858 );
mnot \mul_19_13_g36777/U$1 ( \1860 , \1859 );
mand \mul_19_13_g22509/U$2 ( \1861 , \1847 , \1860 );
mnot \mul_19_13_g22509/U$4 ( \1862 , \1847 );
mand \mul_19_13_g22509/U$3 ( \1863 , \1862 , \1859 );
mnor \mul_19_13_g22509/U$1 ( \1864 , \1861 , \1863 );
mxnor \g37114/U$1_r1 ( \1865 , \1830 , \1864 );
mxor \mul_19_13_g23046/U$1_r1 ( \1866 , \1795 , \1865 );
mxor \g37116/U$1 ( \1867 , \1806 , \1812 );
mxnor \g37116/U$1_r1 ( \1868 , \1867 , \1819 );
mxor \mul_19_13_g22908/U$1 ( \1869 , \b[4] , \c[5] );
mand \g37068/U$2 ( \1870 , \1675 , \1869 );
mand \mul_19_13_g23075/U$1 ( \1871 , \1678 , \1814 );
mnor \g37068/U$1 ( \1872 , \1870 , \1871 );
mnot \mul_19_13_g22534/U$3 ( \1873 , \1728 );
mnot \mul_19_13_g22534/U$4 ( \1874 , \1717 );
mand \mul_19_13_g22534/U$2 ( \1875 , \1873 , \1874 );
mand \mul_19_13_g22534/U$5 ( \1876 , \1728 , \1717 );
mnor \mul_19_13_g22534/U$1 ( \1877 , \1875 , \1876 );
mxor \mul_19_13_g22393/U$4 ( \1878 , \1872 , \1877 );
mnand \mul_19_13_g22675/U$1 ( \1879 , \1773 , \b[0] );
mxor \g36592/U$1 ( \1880 , \c[1] , \b[7] );
mand \g37110/U$2 ( \1881 , \1756 , \1880 );
mand \g37110/U$3 ( \1882 , \1757 , \c[0] );
mnor \g37110/U$1 ( \1883 , \1881 , \1882 );
mxor \mul_19_13_g22489/U$4 ( \1884 , \1879 , \1883 );
mxor \mul_19_13_g22937/U$1 ( \1885 , \b[1] , \c[7] );
mand \mul_19_13_g22623/U$2 ( \1886 , \1782 , \1885 );
mand \mul_19_13_g22623/U$3 ( \1887 , \1747 , \1780 );
mnor \mul_19_13_g22623/U$1 ( \1888 , \1886 , \1887 );
mand \mul_19_13_g22489/U$3 ( \1889 , \1884 , \1888 );
mand \mul_19_13_g22489/U$5 ( \1890 , \1879 , \1883 );
mor \mul_19_13_g22489/U$2 ( \1891 , \1889 , \1890 );
mand \mul_19_13_g22393/U$3 ( \1892 , \1878 , \1891 );
mand \mul_19_13_g22393/U$5 ( \1893 , \1872 , \1877 );
mor \mul_19_13_g22393/U$2 ( \1894 , \1892 , \1893 );
mxor \mul_19_13_g22328/U$4 ( \1895 , \1868 , \1894 );
mxor \mul_19_13_g22409/U$1 ( \1896 , \1729 , \1789 );
mxor \mul_19_13_g22409/U$1_r1 ( \1897 , \1896 , \1792 );
mand \mul_19_13_g22328/U$3 ( \1898 , \1895 , \1897 );
mand \mul_19_13_g22328/U$5 ( \1899 , \1868 , \1894 );
mor \mul_19_13_g22328/U$2 ( \1900 , \1898 , \1899 );
mnand \mul_19_13_g36976/U$1 ( \1901 , \1866 , \1900 );
mxor \mul_19_13_g22328/U$1 ( \1902 , \1868 , \1894 );
mxor \mul_19_13_g22328/U$1_r1 ( \1903 , \1902 , \1897 );
mnot \mul_19_13_g22535/U$3 ( \1904 , \1761 );
mnot \mul_19_13_g22535/U$4 ( \1905 , \1787 );
mor \mul_19_13_g22535/U$2 ( \1906 , \1904 , \1905 );
mnot \mul_19_13_g22551/U$2 ( \1907 , \1787 );
mnand \mul_19_13_g22551/U$1 ( \1908 , \1907 , \1762 );
mnand \mul_19_13_g22535/U$1 ( \1909 , \1906 , \1908 );
mxor \mul_19_13_g23058/U$1 ( \1910 , \1909 , \1776 );
mnot \mul_19_13_g23052/U$2 ( \1911 , \1910 );
mxor \g36593/U$1 ( \1912 , \c[1] , \b[6] );
mnot \mul_19_13_g22686/U$3 ( \1913 , \1912 );
mnot \mul_19_13_g22686/U$4 ( \1914 , \1756 );
mor \mul_19_13_g22686/U$2 ( \1915 , \1913 , \1914 );
mnand \mul_19_13_g22717/U$1 ( \1916 , \1880 , \c[0] );
mnand \mul_19_13_g22686/U$1 ( \1917 , \1915 , \1916 );
mor \mul_19_13_g22820/U$2 ( \1918 , \b[0] , \c[6] );
mnand \mul_19_13_g22820/U$1 ( \1919 , \1918 , \c[5] );
mnand \mul_19_13_g22954/U$1 ( \1920 , \b[0] , \c[6] );
mand \mul_19_13_g22797/U$1 ( \1921 , \1919 , \1920 , \c[7] );
mnand \mul_19_13_g22592/U$1 ( \1922 , \1917 , \1921 );
mxor \mul_19_13_g22919/U$1 ( \1923 , \b[3] , \c[5] );
mnot \mul_19_13_g22642/U$3 ( \1924 , \1923 );
mnot \mul_19_13_g22723/U$2 ( \1925 , \1672 );
mnor \mul_19_13_g22723/U$1 ( \1926 , \1925 , \1674 );
mnot \mul_19_13_g22642/U$4 ( \1927 , \1926 );
mor \mul_19_13_g22642/U$2 ( \1928 , \1924 , \1927 );
mnand \mul_19_13_g22718/U$1 ( \1929 , \1678 , \1869 );
mnand \mul_19_13_g22642/U$1 ( \1930 , \1928 , \1929 );
mnot \mul_19_13_g22641/U$1 ( \1931 , \1930 );
mnand \mul_19_13_g22513/U$1 ( \1932 , \1922 , \1931 );
mxor \mul_19_13_g22903/U$1 ( \1933 , \b[5] , \c[3] );
mnot \mul_19_13_g22659/U$3 ( \1934 , \1933 );
mnot \mul_19_13_g22659/U$4 ( \1935 , \1705 );
mor \mul_19_13_g22659/U$2 ( \1936 , \1934 , \1935 );
mnand \mul_19_13_g22724/U$1 ( \1937 , \1708 , \1719 );
mnand \mul_19_13_g22659/U$1 ( \1938 , \1936 , \1937 );
mand \mul_19_13_g22441/U$2 ( \1939 , \1932 , \1938 );
mnot \mul_19_13_g22544/U$1 ( \1940 , \1922 );
mand \g37045/U$1 ( \1941 , \1940 , \1930 );
mnor \mul_19_13_g22441/U$1 ( \1942 , \1939 , \1941 );
mnand \mul_19_13_g23052/U$1 ( \1943 , \1911 , \1942 );
mnot \mul_19_13_g22341/U$3 ( \1944 , \1943 );
mxor \mul_19_13_g22393/U$1 ( \1945 , \1872 , \1877 );
mxor \mul_19_13_g22393/U$1_r1 ( \1946 , \1945 , \1891 );
mnot \mul_19_13_g22392/U$1 ( \1947 , \1946 );
mnot \mul_19_13_g22341/U$4 ( \1948 , \1947 );
mor \mul_19_13_g22341/U$2 ( \1949 , \1944 , \1948 );
mnot \mul_19_13_g23048/U$2 ( \1950 , \1942 );
mnand \mul_19_13_g23048/U$1 ( \1951 , \1950 , \1910 );
mnand \mul_19_13_g22341/U$1 ( \1952 , \1949 , \1951 );
mnot \mul_19_13_g22334/U$1 ( \1953 , \1952 );
mnand \mul_19_13_g22314/U$1 ( \1954 , \1903 , \1953 );
mxor \mul_19_13_g22489/U$1 ( \1955 , \1879 , \1883 );
mxor \mul_19_13_g22489/U$1_r1 ( \1956 , \1955 , \1888 );
mnot \mul_19_13_g22486/U$1 ( \1957 , \1956 );
mnot \mul_19_13_g22429/U$3 ( \1958 , \1957 );
mxor \mul_19_13_g22904/U$1 ( \1959 , \b[4] , \c[3] );
mnot \mul_19_13_g22664/U$3 ( \1960 , \1959 );
mnot \mul_19_13_g22664/U$4 ( \1961 , \1705 );
mor \mul_19_13_g22664/U$2 ( \1962 , \1960 , \1961 );
mnand \mul_19_13_g22742/U$1 ( \1963 , \1708 , \1933 );
mnand \mul_19_13_g22664/U$1 ( \1964 , \1962 , \1963 );
mxor \mul_19_13_g22920/U$1 ( \1965 , \b[2] , \c[5] );
mnot \mul_19_13_g22648/U$3 ( \1966 , \1965 );
mnot \mul_19_13_g22648/U$4 ( \1967 , \1926 );
mor \mul_19_13_g22648/U$2 ( \1968 , \1966 , \1967 );
mnand \mul_19_13_g22756/U$1 ( \1969 , \1678 , \1923 );
mnand \mul_19_13_g22648/U$1 ( \1970 , \1968 , \1969 );
mor \mul_19_13_g22494/U$2 ( \1971 , \1964 , \1970 );
mxor \mul_19_13_g22943/U$1 ( \1972 , \b[0] , \c[7] );
mnot \mul_19_13_g22628/U$3 ( \1973 , \1972 );
mnot \mul_19_13_g22628/U$4 ( \1974 , \1743 );
mor \mul_19_13_g22628/U$2 ( \1975 , \1973 , \1974 );
mnand \mul_19_13_g22725/U$1 ( \1976 , \1747 , \1885 );
mnand \mul_19_13_g22628/U$1 ( \1977 , \1975 , \1976 );
mnand \mul_19_13_g22494/U$1 ( \1978 , \1971 , \1977 );
mnand \mul_19_13_g22556/U$1 ( \1979 , \1964 , \1970 );
mnand \mul_19_13_g22473/U$1 ( \1980 , \1978 , \1979 );
mnot \mul_19_13_g22456/U$1 ( \1981 , \1980 );
mnot \mul_19_13_g22429/U$4 ( \1982 , \1981 );
mor \mul_19_13_g22429/U$2 ( \1983 , \1958 , \1982 );
mnand \mul_19_13_g22431/U$1 ( \1984 , \1980 , \1956 );
mnand \mul_19_13_g22429/U$1 ( \1985 , \1983 , \1984 );
mnot \mul_19_13_g22504/U$3 ( \1986 , \1931 );
mnot \mul_19_13_g22504/U$4 ( \1987 , \1940 );
mor \mul_19_13_g22504/U$2 ( \1988 , \1986 , \1987 );
mor \mul_19_13_g22504/U$5 ( \1989 , \1940 , \1931 );
mnand \mul_19_13_g22504/U$1 ( \1990 , \1988 , \1989 );
mnot \mul_19_13_g22658/U$1 ( \1991 , \1938 );
mand \mul_19_13_g22442/U$2 ( \1992 , \1990 , \1991 );
mnot \mul_19_13_g22442/U$4 ( \1993 , \1990 );
mand \mul_19_13_g22442/U$3 ( \1994 , \1993 , \1938 );
mnor \mul_19_13_g22442/U$1 ( \1995 , \1992 , \1994 );
mand \mul_19_13_g22396/U$2 ( \1996 , \1985 , \1995 );
mnot \mul_19_13_g22396/U$4 ( \1997 , \1985 );
mnot \mul_19_13_g22422/U$1 ( \1998 , \1995 );
mand \mul_19_13_g22396/U$3 ( \1999 , \1997 , \1998 );
mnor \mul_19_13_g22396/U$1 ( \2000 , \1996 , \1999 );
mxnor \g36585/U$1 ( \2001 , \1917 , \1921 );
mxor \mul_19_13_g22917/U$1 ( \2002 , \b[3] , \c[3] );
mnot \mul_19_13_g22661/U$3 ( \2003 , \2002 );
mnot \mul_19_13_g22661/U$4 ( \2004 , \1705 );
mor \mul_19_13_g22661/U$2 ( \2005 , \2003 , \2004 );
mnand \mul_19_13_g22730/U$1 ( \2006 , \1725 , \1959 );
mnand \mul_19_13_g22661/U$1 ( \2007 , \2005 , \2006 );
mxor \mul_19_13_g22900/U$1 ( \2008 , \b[5] , \c[1] );
mnot \mul_19_13_g22688/U$3 ( \2009 , \2008 );
mnot \mul_19_13_g22688/U$4 ( \2010 , \1756 );
mor \mul_19_13_g22688/U$2 ( \2011 , \2009 , \2010 );
mnand \mul_19_13_g22734/U$1 ( \2012 , \1912 , \c[0] );
mnand \mul_19_13_g22688/U$1 ( \2013 , \2011 , \2012 );
mnot \mul_19_13_g22587/U$2 ( \2014 , \2013 );
mnand \mul_19_13_g22783/U$1 ( \2015 , \1742 , \b[0] );
mnand \mul_19_13_g22587/U$1 ( \2016 , \2014 , \2015 );
mand \mul_19_13_g22497/U$2 ( \2017 , \2007 , \2016 );
mnot \mul_19_13_g22586/U$2 ( \2018 , \2013 );
mnor \mul_19_13_g22586/U$1 ( \2019 , \2018 , \2015 );
mnor \mul_19_13_g22497/U$1 ( \2020 , \2017 , \2019 );
mxor \mul_19_13_g22388/U$4 ( \2021 , \2001 , \2020 );
mxor \mul_19_13_g23065/U$1 ( \2022 , \1977 , \1970 );
mxnor \mul_19_13_g23065/U$1_r1 ( \2023 , \2022 , \1964 );
mand \mul_19_13_g22388/U$3 ( \2024 , \2021 , \2023 );
mand \mul_19_13_g22388/U$5 ( \2025 , \2001 , \2020 );
mor \mul_19_13_g22388/U$2 ( \2026 , \2024 , \2025 );
mnand \mul_19_13_g22337/U$1 ( \2027 , \2000 , \2026 );
mnot \mul_19_13_g22315/U$2 ( \2028 , \2027 );
mnot \mul_19_13_g22395/U$3 ( \2029 , \1942 );
mnot \mul_19_13_g22395/U$4 ( \2030 , \1910 );
mor \mul_19_13_g22395/U$2 ( \2031 , \2029 , \2030 );
mor \mul_19_13_g22395/U$5 ( \2032 , \1942 , \1910 );
mnand \mul_19_13_g22395/U$1 ( \2033 , \2031 , \2032 );
mnot \mul_19_13_g22373/U$1 ( \2034 , \2033 );
mnot \mul_19_13_g22352/U$3 ( \2035 , \2034 );
mnot \mul_19_13_g22352/U$4 ( \2036 , \1947 );
mor \mul_19_13_g22352/U$2 ( \2037 , \2035 , \2036 );
mnand \mul_19_13_g22354/U$1 ( \2038 , \1946 , \2033 );
mnand \mul_19_13_g22352/U$1 ( \2039 , \2037 , \2038 );
mnot \mul_19_13_g22367/U$3 ( \2040 , \1957 );
mnot \mul_19_13_g22367/U$4 ( \2041 , \1998 );
mor \mul_19_13_g22367/U$2 ( \2042 , \2040 , \2041 );
mnot \g37104/U$3 ( \2043 , \1995 );
mnot \g37104/U$4 ( \2044 , \1956 );
mor \g37104/U$2 ( \2045 , \2043 , \2044 );
mnand \g37104/U$1 ( \2046 , \2045 , \1980 );
mnand \mul_19_13_g22367/U$1 ( \2047 , \2042 , \2046 );
mnor \mul_19_13_g22325/U$1 ( \2048 , \2039 , \2047 );
mnor \mul_19_13_g22315/U$1 ( \2049 , \2028 , \2048 );
mand \mul_19_13_g23021/U$1 ( \2050 , \1901 , \1954 , \2049 );
mnot \mul_19_13_g22640/U$3 ( \2051 , \1679 );
mbuf \mul_19_13_g22721/U$1 ( \2052 , \1675 );
mnot \mul_19_13_g22640/U$4 ( \2053 , \2052 );
mor \mul_19_13_g22640/U$2 ( \2054 , \2051 , \2053 );
mxor \mul_19_13_g22885/U$1 ( \2055 , \b[8] , \c[5] );
mnand \mul_19_13_g22712/U$1 ( \2056 , \1678 , \2055 );
mnand \mul_19_13_g22640/U$1 ( \2057 , \2054 , \2056 );
mand \mul_19_13_g22527/U$2 ( \2058 , \1698 , \1711 );
mxor \mul_19_13_g22412/U$1 ( \2059 , \2057 , \2058 );
mnot \mul_19_13_g22522/U$3 ( \2060 , \1843 );
mnot \mul_19_13_g22522/U$4 ( \2061 , \1859 );
mor \mul_19_13_g22522/U$2 ( \2062 , \2060 , \2061 );
mnand \mul_19_13_g22522/U$1 ( \2063 , \2062 , \1836 );
mnot \g36776/U$2 ( \2064 , \1859 );
mnand \g36776/U$1 ( \2065 , \2064 , \1842 );
mnand \mul_19_13_g22498/U$1 ( \2066 , \2063 , \2065 );
mxor \mul_19_13_g22412/U$1_r1 ( \2067 , \2059 , \2066 );
mnot \mul_19_13_g22384/U$3 ( \2068 , \1822 );
mnot \mul_19_13_g22384/U$4 ( \2069 , \1864 );
mor \mul_19_13_g22384/U$2 ( \2070 , \2068 , \2069 );
mor \mul_19_13_g22406/U$2 ( \2071 , \1864 , \1822 );
mnand \mul_19_13_g22406/U$1 ( \2072 , \2071 , \1829 );
mnand \mul_19_13_g22384/U$1 ( \2073 , \2070 , \2072 );
mxor \mul_19_13_g22310/U$1 ( \2074 , \2067 , \2073 );
mxor \mul_19_13_g36691/U$1 ( \2075 , \c[12] , \c[11] );
mand \mul_19_13_g23027/U$1 ( \2076 , \2075 , \b[0] );
mnot \mul_19_13_g22624/U$3 ( \2077 , \1834 );
mnot \mul_19_13_g22624/U$4 ( \2078 , \1782 );
mor \mul_19_13_g22624/U$2 ( \2079 , \2077 , \2078 );
mxor \mul_19_13_g22899/U$1 ( \2080 , \b[6] , \c[7] );
mnand \mul_19_13_g22744/U$1 ( \2081 , \1742 , \2080 );
mnand \mul_19_13_g22624/U$1 ( \2082 , \2079 , \2081 );
mxor \mul_19_13_g22454/U$1 ( \2083 , \2076 , \2082 );
mnot \mul_19_13_g22655/U$3 ( \2084 , \1709 );
mnot \mul_19_13_g22655/U$4 ( \2085 , \1722 );
mor \mul_19_13_g22655/U$2 ( \2086 , \2084 , \2085 );
mxor \mul_19_13_g22856/U$1 ( \2087 , \b[10] , \c[3] );
mnand \mul_19_13_g22743/U$1 ( \2088 , \1725 , \2087 );
mnand \mul_19_13_g22655/U$1 ( \2089 , \2086 , \2088 );
mxor \mul_19_13_g22454/U$1_r1 ( \2090 , \2083 , \2089 );
mnot \g37108/U$3 ( \2091 , \1851 );
mnot \g37108/U$4 ( \2092 , \1857 );
mor \g37108/U$2 ( \2093 , \2091 , \2092 );
mnot \mul_19_13_g37172/U$2 ( \2094 , \c[9] );
mxor \mul_19_13_g37172/U$1 ( \2095 , \b[4] , \2094 );
mnot \mul_19_13_g22672/U$2 ( \2096 , \2095 );
mnand \mul_19_13_g22672/U$1 ( \2097 , \2096 , \1773 );
mnand \g37108/U$1 ( \2098 , \2093 , \2097 );
mnot \mul_19_13_g22704/U$3 ( \2099 , \1840 );
mnot \mul_19_13_g22704/U$4 ( \2100 , \1756 );
mor \mul_19_13_g22704/U$2 ( \2101 , \2099 , \2100 );
mxor \g36589/U$1 ( \2102 , \c[1] , \b[12] );
mnand \mul_19_13_g22780/U$1 ( \2103 , \2102 , \c[0] );
mnand \mul_19_13_g22704/U$1 ( \2104 , \2101 , \2103 );
mxor \mul_19_13_g22510/U$1 ( \2105 , \2098 , \2104 );
mnot \mul_19_13_g22619/U$3 ( \2106 , \1690 );
mnor \mul_19_13_g22812/U$1 ( \2107 , \1689 , \1684 );
mnot \mul_19_13_g22619/U$4 ( \2108 , \2107 );
mor \mul_19_13_g22619/U$2 ( \2109 , \2106 , \2108 );
mxor \mul_19_13_g22940/U$1 ( \2110 , \b[2] , \c[11] );
mnand \mul_19_13_g22748/U$1 ( \2111 , \1689 , \2110 );
mnand \mul_19_13_g22619/U$1 ( \2112 , \2109 , \2111 );
mxor \mul_19_13_g36765/U$1 ( \2113 , \2105 , \2112 );
mxor \mul_19_13_g22350/U$1 ( \2114 , \2090 , \2113 );
mnot \mul_19_13_g22550/U$2 ( \2115 , \1681 );
mnand \mul_19_13_g22550/U$1 ( \2116 , \2115 , \1693 );
mnot \mul_19_13_g22472/U$3 ( \2117 , \2116 );
mnot \mul_19_13_g22472/U$4 ( \2118 , \1712 );
mor \mul_19_13_g22472/U$2 ( \2119 , \2117 , \2118 );
mnand \mul_19_13_g22557/U$1 ( \2120 , \1681 , \1692 );
mnand \mul_19_13_g22472/U$1 ( \2121 , \2119 , \2120 );
mxor \mul_19_13_g22350/U$1_r1 ( \2122 , \2114 , \2121 );
mxor \mul_19_13_g22310/U$1_r1 ( \2123 , \2074 , \2122 );
mnor \mul_19_13_g22360/U$1 ( \2124 , \1794 , \1713 );
mor \mul_19_13_g22332/U$2 ( \2125 , \2124 , \1865 );
mnand \mul_19_13_g22365/U$1 ( \2126 , \1794 , \1713 );
mnand \mul_19_13_g22332/U$1 ( \2127 , \2125 , \2126 );
mnor \mul_19_13_g22292/U$1 ( \2128 , \2123 , \2127 );
mnot \mul_19_13_g22291/U$1 ( \2129 , \2128 );
mxor \mul_19_13_g22388/U$1 ( \2130 , \2001 , \2020 );
mxor \mul_19_13_g22388/U$1_r1 ( \2131 , \2130 , \2023 );
mxor \mul_19_13_g22507/U$1 ( \2132 , \2015 , \2013 );
mxnor \mul_19_13_g22507/U$1_r1 ( \2133 , \2132 , \2007 );
mnand \mul_19_13_g22961/U$1 ( \2134 , \b[0] , \c[4] );
mor \mul_19_13_g22821/U$2 ( \2135 , \b[0] , \c[4] );
mnand \mul_19_13_g22821/U$1 ( \2136 , \2135 , \c[3] );
mnand \mul_19_13_g22795/U$1 ( \2137 , \c[5] , \2134 , \2136 );
mnot \mul_19_13_g23071/U$2 ( \2138 , \2137 );
mxor \mul_19_13_g22902/U$1 ( \2139 , \b[4] , \c[1] );
mnot \mul_19_13_g22687/U$3 ( \2140 , \2139 );
mnot \mul_19_13_g22687/U$4 ( \2141 , \1756 );
mor \mul_19_13_g22687/U$2 ( \2142 , \2140 , \2141 );
mnand \mul_19_13_g22728/U$1 ( \2143 , \2008 , \c[0] );
mnand \mul_19_13_g22687/U$1 ( \2144 , \2142 , \2143 );
mnand \mul_19_13_g23071/U$1 ( \2145 , \2138 , \2144 );
mxor \mul_19_13_g22931/U$1 ( \2146 , \b[1] , \c[5] );
mnot \mul_19_13_g22647/U$3 ( \2147 , \2146 );
mnot \mul_19_13_g22647/U$4 ( \2148 , \1926 );
mor \mul_19_13_g22647/U$2 ( \2149 , \2147 , \2148 );
mnand \mul_19_13_g22765/U$1 ( \2150 , \1678 , \1965 );
mnand \mul_19_13_g22647/U$1 ( \2151 , \2149 , \2150 );
mnot \mul_19_13_g22646/U$1 ( \2152 , \2151 );
mnand \mul_19_13_g22515/U$1 ( \2153 , \2145 , \2152 );
mand \mul_19_13_g22435/U$2 ( \2154 , \2133 , \2153 );
mnot \mul_19_13_g22543/U$1 ( \2155 , \2145 );
mand \mul_19_13_g23022/U$1 ( \2156 , \2155 , \2151 );
mnor \mul_19_13_g22435/U$1 ( \2157 , \2154 , \2156 );
mnand \mul_19_13_g22364/U$1 ( \2158 , \2131 , \2157 );
mnot \mul_19_13_g22279/U$3 ( \2159 , \2158 );
mnot \mul_19_13_g22597/U$3 ( \2160 , \2146 );
mnot \mul_19_13_g22597/U$4 ( \2161 , \1674 );
mor \mul_19_13_g22597/U$2 ( \2162 , \2160 , \2161 );
mxor \mul_19_13_g22945/U$1 ( \2163 , \b[0] , \c[5] );
mnand \mul_19_13_g22741/U$1 ( \2164 , \1672 , \2163 );
mor \mul_19_13_g22597/U$5 ( \2165 , \2164 , \1674 );
mnand \mul_19_13_g22597/U$1 ( \2166 , \2162 , \2165 );
mxor \mul_19_13_g22916/U$1 ( \2167 , \b[2] , \c[3] );
mnot \mul_19_13_g22665/U$3 ( \2168 , \2167 );
mnot \mul_19_13_g22665/U$4 ( \2169 , \1722 );
mor \mul_19_13_g22665/U$2 ( \2170 , \2168 , \2169 );
mnand \mul_19_13_g22753/U$1 ( \2171 , \1725 , \2002 );
mnand \mul_19_13_g22665/U$1 ( \2172 , \2170 , \2171 );
mxor \mul_19_13_g22426/U$4 ( \2173 , \2166 , \2172 );
mnot \g37292/U$2 ( \2174 , \2144 );
mxor \g37292/U$1 ( \2175 , \2137 , \2174 );
mand \mul_19_13_g22426/U$3 ( \2176 , \2173 , \2175 );
mand \mul_19_13_g22426/U$5 ( \2177 , \2166 , \2172 );
mor \mul_19_13_g22426/U$2 ( \2178 , \2176 , \2177 );
mxor \g36573/U$1 ( \2179 , \2155 , \2152 );
mxnor \g36573/U$1_r1 ( \2180 , \2179 , \2133 );
mxor \mul_19_13_g22308/U$4 ( \2181 , \2178 , \2180 );
mxor \g36598/U$1 ( \2182 , \c[1] , \b[2] );
mand \g37111/U$2 ( \2183 , \1756 , \2182 );
mxor \g36597/U$1 ( \2184 , \c[1] , \b[3] );
mand \g37111/U$3 ( \2185 , \2184 , \c[0] );
mnor \g37111/U$1 ( \2186 , \2183 , \2185 );
mor \mul_19_13_g22822/U$2 ( \2187 , \b[0] , \c[2] );
mnand \mul_19_13_g22822/U$1 ( \2188 , \2187 , \c[1] );
mnand \mul_19_13_g22958/U$1 ( \2189 , \b[0] , \c[2] );
mnand \mul_19_13_g22793/U$1 ( \2190 , \2188 , \2189 , \c[3] );
mnot \mul_19_13_g22792/U$1 ( \2191 , \2190 );
mand \mul_19_13_g22578/U$2 ( \2192 , \2186 , \2191 );
mnot \mul_19_13_g22578/U$4 ( \2193 , \2186 );
mand \mul_19_13_g22578/U$3 ( \2194 , \2193 , \2190 );
mnor \mul_19_13_g22578/U$1 ( \2195 , \2192 , \2194 );
mnot \mul_19_13_g22602/U$3 ( \2196 , \1708 );
mxor \mul_19_13_g22949/U$1 ( \2197 , \b[0] , \c[3] );
mnand \mul_19_13_g22755/U$1 ( \2198 , \1702 , \2197 );
mnot \mul_19_13_g22602/U$4 ( \2199 , \2198 );
mand \mul_19_13_g22602/U$2 ( \2200 , \2196 , \2199 );
mxor \mul_19_13_g22929/U$1 ( \2201 , \b[1] , \c[3] );
mand \mul_19_13_g22602/U$5 ( \2202 , \1708 , \2201 );
mnor \mul_19_13_g22602/U$1 ( \2203 , \2200 , \2202 );
mnand \mul_19_13_g22519/U$1 ( \2204 , \2195 , \2203 );
mnot \g37106/U$3 ( \2205 , \2204 );
mand \mul_19_13_g23028/U$1 ( \2206 , \1725 , \b[0] );
mxor \g36599/U$1 ( \2207 , \c[1] , \b[1] );
mnot \mul_19_13_g22693/U$3 ( \2208 , \2207 );
mnot \mul_19_13_g22693/U$4 ( \2209 , \1756 );
mor \mul_19_13_g22693/U$2 ( \2210 , \2208 , \2209 );
mnand \mul_19_13_g22708/U$1 ( \2211 , \2182 , \c[0] );
mnand \mul_19_13_g22693/U$1 ( \2212 , \2210 , \2211 );
mnor \mul_19_13_g22590/U$1 ( \2213 , \2206 , \2212 );
mxor \mul_19_13_g22950/U$1 ( \2214 , \b[0] , \c[1] );
mnot \mul_19_13_g22697/U$3 ( \2215 , \2214 );
mnot \mul_19_13_g22697/U$4 ( \2216 , \1756 );
mor \mul_19_13_g22697/U$2 ( \2217 , \2215 , \2216 );
mnand \mul_19_13_g22757/U$1 ( \2218 , \2207 , \c[0] );
mnand \mul_19_13_g22697/U$1 ( \2219 , \2217 , \2218 );
mnand \mul_19_13_g22977/U$1 ( \2220 , \b[0] , \c[0] );
mand \mul_19_13_g22815/U$1 ( \2221 , \2220 , \c[1] );
mnand \mul_19_13_g22585/U$1 ( \2222 , \2219 , \2221 );
mor \mul_19_13_g22496/U$2 ( \2223 , \2213 , \2222 );
mnand \mul_19_13_g22591/U$1 ( \2224 , \2212 , \2206 );
mnand \mul_19_13_g22496/U$1 ( \2225 , \2223 , \2224 );
mnot \g37106/U$4 ( \2226 , \2225 );
mor \g37106/U$2 ( \2227 , \2205 , \2226 );
mor \mul_19_13_g23056/U$1 ( \2228 , \2195 , \2203 );
mnand \g37106/U$1 ( \2229 , \2227 , \2228 );
mnand \mul_19_13_g22786/U$1 ( \2230 , \1674 , \b[0] );
mnand \mul_19_13_g22767/U$1 ( \2231 , \1702 , \2201 );
mor \mul_19_13_g22600/U$2 ( \2232 , \2231 , \1725 );
mnand \mul_19_13_g22747/U$1 ( \2233 , \2167 , \1703 );
mnand \mul_19_13_g22600/U$1 ( \2234 , \2232 , \2233 );
mnot \mul_19_13_g22599/U$1 ( \2235 , \2234 );
mxor \mul_19_13_g22503/U$1 ( \2236 , \2230 , \2235 );
mnot \mul_19_13_g22690/U$3 ( \2237 , \2184 );
mnot \mul_19_13_g22690/U$4 ( \2238 , \1756 );
mor \mul_19_13_g22690/U$2 ( \2239 , \2237 , \2238 );
mnand \mul_19_13_g22758/U$1 ( \2240 , \2139 , \c[0] );
mnand \mul_19_13_g22690/U$1 ( \2241 , \2239 , \2240 );
mxnor \mul_19_13_g22503/U$1_r1 ( \2242 , \2236 , \2241 );
mnot \mul_19_13_g23067/U$2 ( \2243 , \2186 );
mnand \mul_19_13_g23067/U$1 ( \2244 , \2243 , \2191 );
mnand \mul_19_13_g22448/U$1 ( \2245 , \2242 , \2244 );
mand \mul_19_13_g22381/U$2 ( \2246 , \2229 , \2245 );
mnor \mul_19_13_g22447/U$1 ( \2247 , \2242 , \2244 );
mnor \mul_19_13_g22381/U$1 ( \2248 , \2246 , \2247 );
mxor \mul_19_13_g22426/U$1 ( \2249 , \2166 , \2172 );
mxor \mul_19_13_g22426/U$1_r1 ( \2250 , \2249 , \2175 );
mnot \mul_19_13_g23060/U$2 ( \2251 , \2235 );
mnot \mul_19_13_g22589/U$2 ( \2252 , \2241 );
mnand \mul_19_13_g22589/U$1 ( \2253 , \2252 , \2230 );
mnand \mul_19_13_g23060/U$1 ( \2254 , \2251 , \2253 );
mnot \mul_19_13_g23070/U$2 ( \2255 , \2230 );
mnand \mul_19_13_g23070/U$1 ( \2256 , \2255 , \2241 );
mnand \mul_19_13_g22533/U$1 ( \2257 , \2254 , \2256 );
mnor \mul_19_13_g22401/U$1 ( \2258 , \2250 , \2257 );
mor \mul_19_13_g22340/U$2 ( \2259 , \2248 , \2258 );
mnand \mul_19_13_g22400/U$1 ( \2260 , \2250 , \2257 );
mnand \mul_19_13_g22340/U$1 ( \2261 , \2259 , \2260 );
mand \mul_19_13_g22308/U$3 ( \2262 , \2181 , \2261 );
mand \mul_19_13_g22308/U$5 ( \2263 , \2178 , \2180 );
mor \mul_19_13_g22308/U$2 ( \2264 , \2262 , \2263 );
mnot \mul_19_13_g22279/U$4 ( \2265 , \2264 );
mor \mul_19_13_g22279/U$2 ( \2266 , \2159 , \2265 );
mnot \mul_19_13_g22386/U$1 ( \2267 , \2131 );
mnot \mul_19_13_g22425/U$1 ( \2268 , \2157 );
mnand \mul_19_13_g22362/U$1 ( \2269 , \2267 , \2268 );
mnand \mul_19_13_g22279/U$1 ( \2270 , \2266 , \2269 );
mbuf \mul_19_13_g22268/U$1 ( \2271 , \2270 );
mnand \mul_19_13_g22252/U$1 ( \2272 , \2050 , \2129 , \2271 );
mnor \mul_19_13_g22289/U$1 ( \2273 , \1866 , \1900 );
mnand \g36565/U$1 ( \2274 , \2129 , \2273 );
mnot \mul_19_13_g22358/U$1 ( \2275 , \2000 );
mnot \mul_19_13_g22387/U$1 ( \2276 , \2026 );
mnand \mul_19_13_g22339/U$1 ( \2277 , \2275 , \2276 );
mor \mul_19_13_g22305/U$2 ( \2278 , \2048 , \2277 );
mnand \mul_19_13_g22324/U$1 ( \2279 , \2039 , \2047 );
mnand \mul_19_13_g22305/U$1 ( \2280 , \2278 , \2279 );
mnor \mul_19_13_g22318/U$1 ( \2281 , \1903 , \1953 );
mnor \mul_19_13_g22293/U$1 ( \2282 , \2280 , \2281 );
mnot \mul_19_13_g22267/U$2 ( \2283 , \2282 );
mnand \g36975/U$1 ( \2284 , \1866 , \1900 );
mbuf \fopt36710/U$1 ( \2285 , \1954 );
mnand \mul_19_13_g22267/U$1 ( \2286 , \2283 , \2284 , \2285 , \2129 );
mand \g37048/U$1 ( \2287 , \2123 , \2127 );
mnot \fopt36956/U$1 ( \2288 , \2287 );
mnand \mul_19_13_g22241/U$1 ( \2289 , \2272 , \2274 , \2286 , \2288 );
mnot \mul_19_13_g22700/U$3 ( \2290 , \2102 );
mnot \mul_19_13_g22700/U$4 ( \2291 , \1756 );
mor \mul_19_13_g22700/U$2 ( \2292 , \2290 , \2291 );
mxor \mul_19_13_g22843/U$1 ( \2293 , \b[13] , \c[1] );
mnand \mul_19_13_g22778/U$1 ( \2294 , \2293 , \c[0] );
mnand \mul_19_13_g22700/U$1 ( \2295 , \2292 , \2294 );
mnot \mul_19_13_g22560/U$3 ( \2296 , \2295 );
mor \mul_19_13_g22817/U$2 ( \2297 , \b[0] , \c[12] );
mnand \mul_19_13_g22817/U$1 ( \2298 , \2297 , \c[11] );
mnand \mul_19_13_g22957/U$1 ( \2299 , \b[0] , \c[12] );
mnand \mul_19_13_g22805/U$1 ( \2300 , \2298 , \2299 , \c[13] );
mnot \mul_19_13_g22560/U$4 ( \2301 , \2300 );
mand \mul_19_13_g22560/U$2 ( \2302 , \2296 , \2301 );
mand \mul_19_13_g22560/U$5 ( \2303 , \2295 , \2300 );
mnor \mul_19_13_g22560/U$1 ( \2304 , \2302 , \2303 );
mxor \mul_19_13_g22454/U$4 ( \2305 , \2076 , \2082 );
mand \mul_19_13_g22454/U$3 ( \2306 , \2305 , \2089 );
mand \mul_19_13_g22454/U$5 ( \2307 , \2076 , \2082 );
mor \mul_19_13_g22454/U$2 ( \2308 , \2306 , \2307 );
mxor \mul_19_13_g22385/U$1 ( \2309 , \2304 , \2308 );
mor \mul_19_13_g23057/U$1 ( \2310 , \2098 , \2104 );
mand \mul_19_13_g22452/U$2 ( \2311 , \2310 , \2112 );
mand \mul_19_13_g22510/U$2 ( \2312 , \2098 , \2104 );
mnor \mul_19_13_g22452/U$1 ( \2313 , \2311 , \2312 );
mnot \mul_19_13_g22443/U$1 ( \2314 , \2313 );
mxor \mul_19_13_g22385/U$1_r1 ( \2315 , \2309 , \2314 );
mnot \mul_19_13_g22329/U$3 ( \2316 , \2315 );
mxor \mul_19_13_g22350/U$4 ( \2317 , \2090 , \2113 );
mand \mul_19_13_g22350/U$3 ( \2318 , \2317 , \2121 );
mand \mul_19_13_g22350/U$5 ( \2319 , \2090 , \2113 );
mor \mul_19_13_g22350/U$2 ( \2320 , \2318 , \2319 );
mnot \mul_19_13_g22329/U$4 ( \2321 , \2320 );
mor \mul_19_13_g22329/U$2 ( \2322 , \2316 , \2321 );
mor \mul_19_13_g22329/U$5 ( \2323 , \2320 , \2315 );
mnand \mul_19_13_g22329/U$1 ( \2324 , \2322 , \2323 );
mnot \mul_19_13_g22653/U$3 ( \2325 , \2055 );
mnot \mul_19_13_g22653/U$4 ( \2326 , \1675 );
mor \mul_19_13_g22653/U$2 ( \2327 , \2325 , \2326 );
mxor \mul_19_13_g22884/U$1 ( \2328 , \b[9] , \c[5] );
mnand \mul_19_13_g22764/U$1 ( \2329 , \1678 , \2328 );
mnand \mul_19_13_g22653/U$1 ( \2330 , \2327 , \2329 );
mnot \mul_19_13_g22620/U$3 ( \2331 , \2110 );
mnot \mul_19_13_g22620/U$4 ( \2332 , \1686 );
mor \mul_19_13_g22620/U$2 ( \2333 , \2331 , \2332 );
mxor \mul_19_13_g22939/U$1 ( \2334 , \b[3] , \c[11] );
mnand \mul_19_13_g22766/U$1 ( \2335 , \1689 , \2334 );
mnand \mul_19_13_g22620/U$1 ( \2336 , \2333 , \2335 );
mxor \mul_19_13_g22484/U$1 ( \2337 , \2330 , \2336 );
mxor \mul_19_13_g22913/U$1 ( \2338 , \b[0] , \c[13] );
mnot \mul_19_13_g22609/U$3 ( \2339 , \2338 );
mxnor \mul_19_13_g37188/U$1 ( \2340 , \c[13] , \c[12] );
mnor \mul_19_13_g37241/U$1 ( \2341 , \2340 , \2075 );
mnot \mul_19_13_g22609/U$4 ( \2342 , \2341 );
mor \mul_19_13_g22609/U$2 ( \2343 , \2339 , \2342 );
mxor \mul_19_13_g22942/U$1 ( \2344 , \b[1] , \c[13] );
mnand \mul_19_13_g22713/U$1 ( \2345 , \2075 , \2344 );
mnand \mul_19_13_g22609/U$1 ( \2346 , \2343 , \2345 );
mxor \mul_19_13_g22484/U$1_r1 ( \2347 , \2337 , \2346 );
mnot \mul_19_13_g22483/U$1 ( \2348 , \2347 );
mnot \mul_19_13_g22428/U$3 ( \2349 , \2348 );
mnot \mul_19_13_g22570/U$3 ( \2350 , \1852 );
mnot \mul_19_13_g22570/U$4 ( \2351 , \2095 );
mand \mul_19_13_g22570/U$2 ( \2352 , \2350 , \2351 );
mxor \mul_19_13_g37174/U$1 ( \2353 , \b[5] , \c[9] );
mand \mul_19_13_g22570/U$5 ( \2354 , \1802 , \2353 );
mnor \mul_19_13_g22570/U$1 ( \2355 , \2352 , \2354 );
mnot \mul_19_13_g22569/U$1 ( \2356 , \2355 );
mnot \mul_19_13_g22524/U$3 ( \2357 , \2356 );
mnot \mul_19_13_g22634/U$3 ( \2358 , \2080 );
mnot \mul_19_13_g22634/U$4 ( \2359 , \1743 );
mor \mul_19_13_g22634/U$2 ( \2360 , \2358 , \2359 );
mxor \mul_19_13_g22898/U$1 ( \2361 , \b[7] , \c[7] );
mnand \mul_19_13_g22754/U$1 ( \2362 , \1747 , \2361 );
mnand \mul_19_13_g22634/U$1 ( \2363 , \2360 , \2362 );
mnot \mul_19_13_g22633/U$1 ( \2364 , \2363 );
mnot \mul_19_13_g22524/U$4 ( \2365 , \2364 );
mor \mul_19_13_g22524/U$2 ( \2366 , \2357 , \2365 );
mnand \mul_19_13_g22530/U$1 ( \2367 , \2355 , \2363 );
mnand \mul_19_13_g22524/U$1 ( \2368 , \2366 , \2367 );
mnot \mul_19_13_g22657/U$3 ( \2369 , \2087 );
mbuf \mul_19_13_g22759/U$1 ( \2370 , \1705 );
mnot \mul_19_13_g22657/U$4 ( \2371 , \2370 );
mor \mul_19_13_g22657/U$2 ( \2372 , \2369 , \2371 );
mxor \mul_19_13_g22857/U$1 ( \2373 , \b[11] , \c[3] );
mnand \mul_19_13_g22750/U$1 ( \2374 , \1708 , \2373 );
mnand \mul_19_13_g22657/U$1 ( \2375 , \2372 , \2374 );
mxnor \mul_19_13_g23064/U$1 ( \2376 , \2368 , \2375 );
mnot \mul_19_13_g22457/U$1 ( \2377 , \2376 );
mnot \mul_19_13_g22428/U$4 ( \2378 , \2377 );
mor \mul_19_13_g22428/U$2 ( \2379 , \2349 , \2378 );
mnand \mul_19_13_g22430/U$1 ( \2380 , \2376 , \2347 );
mnand \mul_19_13_g22428/U$1 ( \2381 , \2379 , \2380 );
mxor \mul_19_13_g22412/U$4 ( \2382 , \2057 , \2058 );
mand \mul_19_13_g22412/U$3 ( \2383 , \2382 , \2066 );
mand \mul_19_13_g22412/U$5 ( \2384 , \2057 , \2058 );
mor \mul_19_13_g22412/U$2 ( \2385 , \2383 , \2384 );
mnot \mul_19_13_g22411/U$1 ( \2386 , \2385 );
mand \mul_19_13_g22375/U$2 ( \2387 , \2381 , \2386 );
mnot \mul_19_13_g22375/U$4 ( \2388 , \2381 );
mand \mul_19_13_g22375/U$3 ( \2389 , \2388 , \2385 );
mnor \mul_19_13_g22375/U$1 ( \2390 , \2387 , \2389 );
mand \mul_19_13_g22311/U$2 ( \2391 , \2324 , \2390 );
mnot \mul_19_13_g22311/U$4 ( \2392 , \2324 );
mnot \mul_19_13_g22346/U$1 ( \2393 , \2390 );
mand \mul_19_13_g22311/U$3 ( \2394 , \2392 , \2393 );
mnor \mul_19_13_g22311/U$1 ( \2395 , \2391 , \2394 );
mnot \mul_19_13_g23037/U$2 ( \2396 , \2395 );
mxor \mul_19_13_g22310/U$4 ( \2397 , \2067 , \2073 );
mand \mul_19_13_g22310/U$3 ( \2398 , \2397 , \2122 );
mand \mul_19_13_g22310/U$5 ( \2399 , \2067 , \2073 );
mor \mul_19_13_g22310/U$2 ( \2400 , \2398 , \2399 );
mnand \mul_19_13_g23037/U$1 ( \2401 , \2396 , \2400 );
mnot \mul_19_13_g22274/U$2 ( \2402 , \2400 );
mnand \mul_19_13_g22274/U$1 ( \2403 , \2402 , \2395 );
mnand \mul_19_13_g22263/U$1 ( \2404 , \2401 , \2403 );
mnot \mul_19_13_g22262/U$1 ( \2405 , \2404 );
mand \mul_19_13_g22236/U$2 ( \2406 , \2289 , \2405 );
mnot \mul_19_13_g22236/U$4 ( \2407 , \2289 );
mand \mul_19_13_g22236/U$3 ( \2408 , \2407 , \2404 );
mnor \mul_19_13_g22236/U$1 ( \2409 , \2406 , \2408 );
mxor \mul_6_11_g6500/U$1 ( \2410 , \155 , \202 );
mxor \mul_6_11_g6500/U$1_r1 ( \2411 , \2410 , \344 );
mnot \g4816/U$1 ( \2412 , \2411 );
mnot \g4815/U$1 ( \2413 , \2412 );
mnand \g4753/U$1 ( \2414 , \2409 , \2413 );
mor \g4759/U$1 ( \2415 , \a[13] , \d[13] );
mnot \g4651/U$3 ( \2416 , \2415 );
mnot \g4651/U$4 ( \2417 , \648 );
mor \g4651/U$2 ( \2418 , \2416 , \2417 );
mor \g4757/U$1 ( \2419 , \a[13] , \b[13] );
mnand \g4687/U$1 ( \2420 , \667 , \2419 );
mnand \g4651/U$1 ( \2421 , \2418 , \2420 );
mand \g4761/U$1 ( \2422 , \b[13] , \c[13] );
mnot \g4585/U$3 ( \2423 , \2422 );
mnot \g4585/U$4 ( \2424 , \922 );
mor \g4585/U$2 ( \2425 , \2423 , \2424 );
mxor \g4725/U$1 ( \2426 , \c[13] , \d[13] );
mand \g4612/U$2 ( \2427 , \697 , \2426 );
mnot \add_17_12_g6763/U$2 ( \2428 , \757 );
mnand \add_17_12_g6763/U$1 ( \2429 , \2428 , \781 );
mnot \add_17_12_g6689/U$3 ( \2430 , \2429 );
mor \add_17_12_g6696/U$2 ( \2431 , \777 , \758 );
mnot \add_17_12_g6703/U$2 ( \2432 , \758 );
mnand \add_17_12_g6703/U$1 ( \2433 , \2432 , \747 , \754 );
mnand \add_17_12_g6696/U$1 ( \2434 , \2431 , \2433 , \779 );
mnot \add_17_12_g6689/U$4 ( \2435 , \2434 );
mor \add_17_12_g6689/U$2 ( \2436 , \2430 , \2435 );
mor \add_17_12_g6689/U$5 ( \2437 , \2434 , \2429 );
mnand \add_17_12_g6689/U$1 ( \2438 , \2436 , \2437 );
mnot \g4621/U$3 ( \2439 , \2438 );
mnot \g4621/U$4 ( \2440 , \707 );
mor \g4621/U$2 ( \2441 , \2439 , \2440 );
mnot \add_16_12_g6763/U$2 ( \2442 , \842 );
mnand \add_16_12_g6763/U$1 ( \2443 , \2442 , \866 );
mnot \add_16_12_g6689/U$3 ( \2444 , \2443 );
mor \add_16_12_g6696/U$2 ( \2445 , \862 , \843 );
mnot \add_16_12_g6703/U$2 ( \2446 , \843 );
mnand \add_16_12_g6703/U$1 ( \2447 , \2446 , \832 , \839 );
mnand \add_16_12_g6696/U$1 ( \2448 , \2445 , \2447 , \864 );
mnot \add_16_12_g6689/U$4 ( \2449 , \2448 );
mor \add_16_12_g6689/U$2 ( \2450 , \2444 , \2449 );
mor \add_16_12_g6689/U$5 ( \2451 , \2448 , \2443 );
mnand \add_16_12_g6689/U$1 ( \2452 , \2450 , \2451 );
mand \g4643/U$2 ( \2453 , \880 , \2452 );
mnot \g4668/U$3 ( \2454 , \d[13] );
mnot \g4668/U$4 ( \2455 , \894 );
mor \g4668/U$2 ( \2456 , \2454 , \2455 );
mand \g4707/U$2 ( \2457 , \885 , \b[13] );
mand \g4707/U$3 ( \2458 , \907 , \c[13] );
mnor \g4707/U$1 ( \2459 , \2457 , \2458 );
mnand \g4668/U$1 ( \2460 , \2456 , \2459 );
mnor \g4643/U$1 ( \2461 , \2453 , \2460 );
mnand \g4621/U$1 ( \2462 , \2441 , \2461 );
mnor \g4612/U$1 ( \2463 , \2427 , \2462 );
mnand \g4585/U$1 ( \2464 , \2425 , \2463 );
mnor \g4582/U$1 ( \2465 , \2421 , \2464 );
mxor \g36943/U$1 ( \2466 , \915 , \916 );
mnot \g4914/U$2 ( \2467 , \705 );
mnor \g4792/U$1 ( \2468 , \907 , \885 );
mnand \g4692/U$1 ( \2469 , \893 , \2468 );
mnor \g4666/U$1 ( \2470 , \879 , \2469 );
mnand \g4914/U$1 ( \2471 , \2467 , \2470 );
mnor \g4629/U$1 ( \2472 , \1666 , \2471 );
mnand \g4599/U$1 ( \2473 , \2412 , \2472 );
mnor \g4588/U$1 ( \2474 , \2473 , \695 );
mand \g4909/U$1 ( \2475 , \2466 , \2474 );
mnand \g4543/U$1 ( \2476 , \2475 , \a[13] );
mnand \g4515/U$1 ( \2477 , \1669 , \2414 , \2465 , \2476 );
mnot \mul_19_13_g22608/U$3 ( \2478 , \2344 );
mnot \mul_19_13_g22608/U$4 ( \2479 , \2341 );
mor \mul_19_13_g22608/U$2 ( \2480 , \2478 , \2479 );
mxor \mul_19_13_g22947/U$1 ( \2481 , \b[2] , \c[13] );
mnand \mul_19_13_g22739/U$1 ( \2482 , \2075 , \2481 );
mnand \mul_19_13_g22608/U$1 ( \2483 , \2480 , \2482 );
mnot \mul_19_13_g23073/U$2 ( \2484 , \2300 );
mnand \mul_19_13_g23073/U$1 ( \2485 , \2484 , \2295 );
mxor \mul_19_13_g22445/U$1 ( \2486 , \2483 , \2485 );
mnot \mul_19_13_g22617/U$3 ( \2487 , \2334 );
mnot \mul_19_13_g22617/U$4 ( \2488 , \2107 );
mor \mul_19_13_g22617/U$2 ( \2489 , \2487 , \2488 );
mxor \mul_19_13_g22933/U$1 ( \2490 , \b[4] , \c[11] );
mnand \mul_19_13_g22735/U$1 ( \2491 , \1689 , \2490 );
mnand \mul_19_13_g22617/U$1 ( \2492 , \2489 , \2491 );
mxor \mul_19_13_g22445/U$1_r1 ( \2493 , \2486 , \2492 );
mnot \mul_19_13_g22420/U$1 ( \2494 , \2493 );
mnot \mul_19_13_g22394/U$3 ( \2495 , \2494 );
mnot \g37107/U$3 ( \2496 , \1773 );
mxor \mul_19_13_g22905/U$1 ( \2497 , \b[6] , \c[9] );
mnot \g37107/U$4 ( \2498 , \2497 );
mor \g37107/U$2 ( \2499 , \2496 , \2498 );
mnand \mul_19_13_g22581/U$1 ( \2500 , \1770 , \2353 );
mnand \g37107/U$1 ( \2501 , \2499 , \2500 );
mnot \mul_19_13_g22631/U$3 ( \2502 , \2361 );
mnot \mul_19_13_g22631/U$4 ( \2503 , \1743 );
mor \mul_19_13_g22631/U$2 ( \2504 , \2502 , \2503 );
mxor \mul_19_13_g22888/U$1 ( \2505 , \b[8] , \c[7] );
mnand \mul_19_13_g22746/U$1 ( \2506 , \1747 , \2505 );
mnand \mul_19_13_g22631/U$1 ( \2507 , \2504 , \2506 );
mxor \mul_19_13_g22463/U$1 ( \2508 , \2501 , \2507 );
mnot \mul_19_13_g22649/U$3 ( \2509 , \2328 );
mnot \mul_19_13_g22649/U$4 ( \2510 , \2052 );
mor \mul_19_13_g22649/U$2 ( \2511 , \2509 , \2510 );
mxor \mul_19_13_g22859/U$1 ( \2512 , \b[10] , \c[5] );
mnand \mul_19_13_g22740/U$1 ( \2513 , \1678 , \2512 );
mnand \mul_19_13_g22649/U$1 ( \2514 , \2511 , \2513 );
mxor \mul_19_13_g22463/U$1_r1 ( \2515 , \2508 , \2514 );
mnot \mul_19_13_g22459/U$1 ( \2516 , \2515 );
mnot \mul_19_13_g22394/U$4 ( \2517 , \2516 );
mor \mul_19_13_g22394/U$2 ( \2518 , \2495 , \2517 );
mnand \mul_19_13_g22398/U$1 ( \2519 , \2493 , \2515 );
mnand \mul_19_13_g22394/U$1 ( \2520 , \2518 , \2519 );
mnot \mul_19_13_g22405/U$3 ( \2521 , \2304 );
mnot \mul_19_13_g22405/U$4 ( \2522 , \2313 );
mor \mul_19_13_g22405/U$2 ( \2523 , \2521 , \2522 );
mnand \mul_19_13_g22405/U$1 ( \2524 , \2523 , \2308 );
mnot \mul_19_13_g22415/U$2 ( \2525 , \2304 );
mnand \mul_19_13_g22415/U$1 ( \2526 , \2525 , \2314 );
mnand \mul_19_13_g22379/U$1 ( \2527 , \2524 , \2526 );
mxnor \mul_19_13_g23045/U$1 ( \2528 , \2520 , \2527 );
mnot \mul_19_13_g22321/U$3 ( \2529 , \2528 );
mxor \mul_19_13_g22484/U$4 ( \2530 , \2330 , \2336 );
mand \mul_19_13_g22484/U$3 ( \2531 , \2530 , \2346 );
mand \mul_19_13_g22484/U$5 ( \2532 , \2330 , \2336 );
mor \mul_19_13_g22484/U$2 ( \2533 , \2531 , \2532 );
mxor \mul_19_13_g22887/U$1 ( \2534 , \c[14] , \c[13] );
mand \mul_19_13_g23023/U$1 ( \2535 , \2534 , \b[0] );
mnot \mul_19_13_g22701/U$3 ( \2536 , \1756 );
mnot \mul_19_13_g22701/U$4 ( \2537 , \2293 );
mor \mul_19_13_g22701/U$2 ( \2538 , \2536 , \2537 );
mxor \mul_19_13_g23076/U$1 ( \2539 , \c[1] , \b[14] );
mnand \mul_19_13_g22779/U$1 ( \2540 , \2539 , \c[0] );
mnand \mul_19_13_g22701/U$1 ( \2541 , \2538 , \2540 );
mxor \mul_19_13_g22485/U$1 ( \2542 , \2535 , \2541 );
mnot \mul_19_13_g22669/U$3 ( \2543 , \2373 );
mnot \mul_19_13_g22669/U$4 ( \2544 , \1705 );
mor \mul_19_13_g22669/U$2 ( \2545 , \2543 , \2544 );
mxor \mul_19_13_g22847/U$1 ( \2546 , \b[12] , \c[3] );
mnand \mul_19_13_g22789/U$1 ( \2547 , \1708 , \2546 );
mnand \mul_19_13_g22669/U$1 ( \2548 , \2545 , \2547 );
mxor \mul_19_13_g22485/U$1_r1 ( \2549 , \2542 , \2548 );
mxor \mul_19_13_g22369/U$1 ( \2550 , \2533 , \2549 );
mor \mul_19_13_g22521/U$2 ( \2551 , \2375 , \2356 );
mnand \mul_19_13_g22521/U$1 ( \2552 , \2551 , \2363 );
mnand \mul_19_13_g22528/U$1 ( \2553 , \2375 , \2356 );
mnand \mul_19_13_g22500/U$1 ( \2554 , \2552 , \2553 );
mxor \mul_19_13_g22369/U$1_r1 ( \2555 , \2550 , \2554 );
mnot \mul_19_13_g22321/U$4 ( \2556 , \2555 );
mand \mul_19_13_g22321/U$2 ( \2557 , \2529 , \2556 );
mand \mul_19_13_g22321/U$5 ( \2558 , \2528 , \2555 );
mnor \mul_19_13_g22321/U$1 ( \2559 , \2557 , \2558 );
mnot \mul_19_13_g22284/U$3 ( \2560 , \2559 );
mnot \mul_19_13_g22357/U$3 ( \2561 , \2347 );
mnot \mul_19_13_g22357/U$4 ( \2562 , \2385 );
mor \mul_19_13_g22357/U$2 ( \2563 , \2561 , \2562 );
mor \mul_19_13_g22366/U$2 ( \2564 , \2385 , \2347 );
mnand \mul_19_13_g22366/U$1 ( \2565 , \2564 , \2377 );
mnand \mul_19_13_g22357/U$1 ( \2566 , \2563 , \2565 );
mnot \mul_19_13_g22284/U$4 ( \2567 , \2566 );
mand \mul_19_13_g22284/U$2 ( \2568 , \2560 , \2567 );
mand \mul_19_13_g22284/U$5 ( \2569 , \2559 , \2566 );
mnor \mul_19_13_g22284/U$1 ( \2570 , \2568 , \2569 );
mnot \mul_19_13_g23035/U$2 ( \2571 , \2570 );
mnot \mul_19_13_g22326/U$3 ( \2572 , \2315 );
mnot \mul_19_13_g22326/U$4 ( \2573 , \2390 );
mor \mul_19_13_g22326/U$2 ( \2574 , \2572 , \2573 );
mnand \mul_19_13_g22326/U$1 ( \2575 , \2574 , \2320 );
mnot \mul_19_13_g23044/U$2 ( \2576 , \2315 );
mnand \mul_19_13_g23044/U$1 ( \2577 , \2576 , \2393 );
mnand \mul_19_13_g22320/U$1 ( \2578 , \2575 , \2577 );
mnand \mul_19_13_g23035/U$1 ( \2579 , \2571 , \2578 );
mnot \mul_19_13_g22258/U$2 ( \2580 , \2578 );
mnand \mul_19_13_g22258/U$1 ( \2581 , \2580 , \2570 );
mnand \mul_19_13_g22248/U$1 ( \2582 , \2579 , \2581 );
mnot \mul_19_13_g22232/U$3 ( \2583 , \2582 );
mand \mul_19_13_g2/U$1 ( \2584 , \2129 , \2403 , \1901 );
mnot \mul_19_13_g22234/U$3 ( \2585 , \2584 );
mnot \g37264/U$2 ( \2586 , \2273 );
mnand \mul_19_13_g22257/U$1 ( \2587 , \2270 , \2049 );
mnot \mul_19_13_g22245/U$3 ( \2588 , \2587 );
mnot \mul_19_13_g22245/U$4 ( \2589 , \2282 );
mor \mul_19_13_g22245/U$2 ( \2590 , \2588 , \2589 );
mnand \mul_19_13_g22245/U$1 ( \2591 , \2590 , \2285 );
mnand \g37264/U$1 ( \2592 , \2586 , \2591 );
mnot \mul_19_13_g22234/U$4 ( \2593 , \2592 );
mor \mul_19_13_g22234/U$2 ( \2594 , \2585 , \2593 );
mnand \mul_19_13_g22264/U$1 ( \2595 , \2287 , \2403 );
mnand \mul_19_13_g22260/U$1 ( \2596 , \2595 , \2401 );
mnot \mul_19_13_g22259/U$1 ( \2597 , \2596 );
mnand \mul_19_13_g22234/U$1 ( \2598 , \2594 , \2597 );
mnot \mul_19_13_g22232/U$4 ( \2599 , \2598 );
mor \mul_19_13_g22232/U$2 ( \2600 , \2583 , \2599 );
mor \mul_19_13_g22232/U$5 ( \2601 , \2582 , \2598 );
mnand \mul_19_13_g22232/U$1 ( \2602 , \2600 , \2601 );
mnand \g4789/U$1 ( \2603 , \2602 , \2413 );
mnot \g4655/U$3 ( \2604 , \686 );
mnot \g4655/U$4 ( \2605 , \648 );
mor \g4655/U$2 ( \2606 , \2604 , \2605 );
mor \g37083/U$2 ( \2607 , \a[14] , \b[14] );
mnand \g37083/U$1 ( \2608 , \2607 , \667 );
mnand \g4655/U$1 ( \2609 , \2606 , \2608 );
mand \g4737/U$1 ( \2610 , \b[14] , \c[14] );
mnot \g4584/U$3 ( \2611 , \2610 );
mnot \g4584/U$4 ( \2612 , \922 );
mor \g4584/U$2 ( \2613 , \2611 , \2612 );
mnot \g4830/U$1 ( \2614 , \696 );
mbuf \g4829/U$1 ( \2615 , \2614 );
mxor \g4734/U$1 ( \2616 , \c[14] , \d[14] );
mand \g4611/U$2 ( \2617 , \2615 , \2616 );
mnot \add_17_12_g6758/U$2 ( \2618 , \785 );
mnor \add_17_12_g6758/U$1 ( \2619 , \2618 , \755 );
mnot \add_17_12_g6688/U$3 ( \2620 , \2619 );
mand \add_17_12_g6699/U$2 ( \2621 , \747 , \754 , \759 );
mnot \add_17_12_g6712/U$2 ( \2622 , \782 );
mnand \add_17_12_g6718/U$1 ( \2623 , \776 , \759 );
mnand \add_17_12_g6712/U$1 ( \2624 , \2622 , \2623 );
mnor \add_17_12_g6699/U$1 ( \2625 , \2621 , \2624 );
mnot \add_17_12_g6688/U$4 ( \2626 , \2625 );
mor \add_17_12_g6688/U$2 ( \2627 , \2620 , \2626 );
mor \add_17_12_g6688/U$5 ( \2628 , \2625 , \2619 );
mnand \add_17_12_g6688/U$1 ( \2629 , \2627 , \2628 );
mnot \g4616/U$3 ( \2630 , \2629 );
mnot \g4616/U$4 ( \2631 , \707 );
mor \g4616/U$2 ( \2632 , \2630 , \2631 );
mnot \add_16_12_g6758/U$2 ( \2633 , \870 );
mnor \add_16_12_g6758/U$1 ( \2634 , \2633 , \840 );
mnot \add_16_12_g6688/U$3 ( \2635 , \2634 );
mand \add_16_12_g6699/U$2 ( \2636 , \832 , \839 , \844 );
mnot \add_16_12_g6712/U$2 ( \2637 , \867 );
mnand \add_16_12_g6718/U$1 ( \2638 , \861 , \844 );
mnand \add_16_12_g6712/U$1 ( \2639 , \2637 , \2638 );
mnor \add_16_12_g6699/U$1 ( \2640 , \2636 , \2639 );
mnot \add_16_12_g6688/U$4 ( \2641 , \2640 );
mor \add_16_12_g6688/U$2 ( \2642 , \2635 , \2641 );
mor \add_16_12_g6688/U$5 ( \2643 , \2640 , \2634 );
mnand \add_16_12_g6688/U$1 ( \2644 , \2642 , \2643 );
mand \g4637/U$2 ( \2645 , \880 , \2644 );
mnot \g4662/U$3 ( \2646 , \d[14] );
mnot \g4662/U$4 ( \2647 , \894 );
mor \g4662/U$2 ( \2648 , \2646 , \2647 );
mand \g4703/U$2 ( \2649 , \885 , \b[14] );
mand \g4703/U$3 ( \2650 , \907 , \c[14] );
mnor \g4703/U$1 ( \2651 , \2649 , \2650 );
mnand \g4662/U$1 ( \2652 , \2648 , \2651 );
mnor \g4637/U$1 ( \2653 , \2645 , \2652 );
mnand \g4616/U$1 ( \2654 , \2632 , \2653 );
mnor \g4611/U$1 ( \2655 , \2617 , \2654 );
mnand \g4584/U$1 ( \2656 , \2613 , \2655 );
mnor \g4568/U$1 ( \2657 , \2609 , \2656 );
mnot \mul_18_12_g22608/U$3 ( \2658 , \1586 );
mnor \mul_18_12_g22808/U$1 ( \2659 , \1582 , \1335 );
mnot \mul_18_12_g22608/U$4 ( \2660 , \2659 );
mor \mul_18_12_g22608/U$2 ( \2661 , \2658 , \2660 );
mxor \mul_18_12_g22947/U$1 ( \2662 , \a[2] , \d[13] );
mnand \mul_18_12_g22739/U$1 ( \2663 , \1335 , \2662 );
mnand \mul_18_12_g22608/U$1 ( \2664 , \2661 , \2663 );
mnot \mul_18_12_g23073/U$2 ( \2665 , \1555 );
mnand \mul_18_12_g23073/U$1 ( \2666 , \2665 , \1550 );
mxor \mul_18_12_g22445/U$1 ( \2667 , \2664 , \2666 );
mnot \mul_18_12_g22617/U$3 ( \2668 , \1592 );
mnot \mul_18_12_g22617/U$4 ( \2669 , \1366 );
mor \mul_18_12_g22617/U$2 ( \2670 , \2668 , \2669 );
mxor \mul_18_12_g22933/U$1 ( \2671 , \a[4] , \d[11] );
mnand \mul_18_12_g22735/U$1 ( \2672 , \947 , \2671 );
mnand \mul_18_12_g22617/U$1 ( \2673 , \2670 , \2672 );
mxor \mul_18_12_g22445/U$1_r1 ( \2674 , \2667 , \2673 );
mnot \fopt36952/U$1 ( \2675 , \2674 );
mnot \mul_18_12_g22394/U$3 ( \2676 , \2675 );
mnot \g37123/U$3 ( \2677 , \1026 );
mnot \g37123/U$4 ( \2678 , \1608 );
mor \g37123/U$2 ( \2679 , \2677 , \2678 );
mxor \mul_18_12_g22905/U$1 ( \2680 , \a[6] , \d[9] );
mnand \mul_18_12_g22674/U$1 ( \2681 , \1029 , \2680 );
mnand \g37123/U$1 ( \2682 , \2679 , \2681 );
mnot \mul_18_12_g22631/U$3 ( \2683 , \1616 );
mnot \mul_18_12_g22631/U$4 ( \2684 , \999 );
mor \mul_18_12_g22631/U$2 ( \2685 , \2683 , \2684 );
mxor \mul_18_12_g22888/U$1 ( \2686 , \a[8] , \d[7] );
mnand \mul_18_12_g22746/U$1 ( \2687 , \1003 , \2686 );
mnand \mul_18_12_g22631/U$1 ( \2688 , \2685 , \2687 );
mxor \mul_18_12_g22463/U$1 ( \2689 , \2682 , \2688 );
mnot \mul_18_12_g22649/U$3 ( \2690 , \1599 );
mnot \mul_18_12_g22649/U$4 ( \2691 , \1312 );
mor \mul_18_12_g22649/U$2 ( \2692 , \2690 , \2691 );
mxor \mul_18_12_g22859/U$1 ( \2693 , \a[10] , \d[5] );
mnand \mul_18_12_g22740/U$1 ( \2694 , \936 , \2693 );
mnand \mul_18_12_g22649/U$1 ( \2695 , \2692 , \2694 );
mxor \mul_18_12_g22463/U$1_r1 ( \2696 , \2689 , \2695 );
mnot \mul_18_12_g22459/U$1 ( \2697 , \2696 );
mnot \mul_18_12_g22394/U$4 ( \2698 , \2697 );
mor \mul_18_12_g22394/U$2 ( \2699 , \2676 , \2698 );
mnand \mul_18_12_g22398/U$1 ( \2700 , \2674 , \2696 );
mnand \mul_18_12_g22394/U$1 ( \2701 , \2699 , \2700 );
mnot \mul_18_12_g22405/U$3 ( \2702 , \1559 );
mnot \mul_18_12_g22405/U$4 ( \2703 , \1568 );
mor \mul_18_12_g22405/U$2 ( \2704 , \2702 , \2703 );
mnand \mul_18_12_g22405/U$1 ( \2705 , \2704 , \1563 );
mnot \mul_18_12_g22415/U$2 ( \2706 , \1559 );
mnand \mul_18_12_g22415/U$1 ( \2707 , \2706 , \1569 );
mnand \mul_18_12_g22379/U$1 ( \2708 , \2705 , \2707 );
mxnor \mul_18_12_g23045/U$1 ( \2709 , \2701 , \2708 );
mnot \mul_18_12_g22321/U$3 ( \2710 , \2709 );
mxor \mul_18_12_g22484/U$4 ( \2711 , \1588 , \1594 );
mand \mul_18_12_g22484/U$3 ( \2712 , \2711 , \1601 );
mand \mul_18_12_g22484/U$5 ( \2713 , \1588 , \1594 );
mor \mul_18_12_g22484/U$2 ( \2714 , \2712 , \2713 );
mxor \mul_18_12_g22887/U$1 ( \2715 , \d[14] , \d[13] );
mand \mul_18_12_g23023/U$1 ( \2716 , \2715 , \a[0] );
mnot \mul_18_12_g22701/U$3 ( \2717 , \1012 );
mnot \mul_18_12_g22701/U$4 ( \2718 , \1548 );
mor \mul_18_12_g22701/U$2 ( \2719 , \2717 , \2718 );
mxor \mul_18_12_g23076/U$1 ( \2720 , \d[1] , \a[14] );
mnand \mul_18_12_g22779/U$1 ( \2721 , \2720 , \d[0] );
mnand \mul_18_12_g22701/U$1 ( \2722 , \2719 , \2721 );
mxor \mul_18_12_g22485/U$1 ( \2723 , \2716 , \2722 );
mnot \mul_18_12_g22669/U$3 ( \2724 , \1627 );
mnot \mul_18_12_g22669/U$4 ( \2725 , \962 );
mor \mul_18_12_g22669/U$2 ( \2726 , \2724 , \2725 );
mxor \mul_18_12_g22847/U$1 ( \2727 , \a[12] , \d[3] );
mnand \mul_18_12_g22789/U$1 ( \2728 , \965 , \2727 );
mnand \mul_18_12_g22669/U$1 ( \2729 , \2726 , \2728 );
mxor \mul_18_12_g22485/U$1_r1 ( \2730 , \2723 , \2729 );
mxor \mul_18_12_g22369/U$1 ( \2731 , \2714 , \2730 );
mnot \fopt36731/U$1 ( \2732 , \1610 );
mnand \mul_18_12_g22528/U$1 ( \2733 , \1629 , \2732 );
mor \mul_18_12_g22521/U$2 ( \2734 , \1629 , \2732 );
mnand \mul_18_12_g22521/U$1 ( \2735 , \2734 , \1618 );
mnand \mul_18_12_g22500/U$1 ( \2736 , \2733 , \2735 );
mxor \mul_18_12_g22369/U$1_r1 ( \2737 , \2731 , \2736 );
mnot \mul_18_12_g22321/U$4 ( \2738 , \2737 );
mand \mul_18_12_g22321/U$2 ( \2739 , \2710 , \2738 );
mand \mul_18_12_g22321/U$5 ( \2740 , \2709 , \2737 );
mnor \mul_18_12_g22321/U$1 ( \2741 , \2739 , \2740 );
mnot \mul_18_12_g22284/U$3 ( \2742 , \2741 );
mnot \mul_18_12_g22357/U$3 ( \2743 , \1602 );
mnot \mul_18_12_g22357/U$4 ( \2744 , \1639 );
mor \mul_18_12_g22357/U$2 ( \2745 , \2743 , \2744 );
mor \mul_18_12_g22366/U$2 ( \2746 , \1639 , \1602 );
mnand \mul_18_12_g22366/U$1 ( \2747 , \2746 , \1631 );
mnand \mul_18_12_g22357/U$1 ( \2748 , \2745 , \2747 );
mnot \mul_18_12_g22284/U$4 ( \2749 , \2748 );
mand \mul_18_12_g22284/U$2 ( \2750 , \2742 , \2749 );
mand \mul_18_12_g22284/U$5 ( \2751 , \2741 , \2748 );
mnor \mul_18_12_g22284/U$1 ( \2752 , \2750 , \2751 );
mnot \mul_18_12_g23035/U$2 ( \2753 , \2752 );
mnot \mul_18_12_g22326/U$3 ( \2754 , \1570 );
mnot \mul_18_12_g22326/U$4 ( \2755 , \1644 );
mor \mul_18_12_g22326/U$2 ( \2756 , \2754 , \2755 );
mnand \mul_18_12_g22326/U$1 ( \2757 , \2756 , \1575 );
mnot \mul_18_12_g23044/U$2 ( \2758 , \1570 );
mnand \mul_18_12_g23044/U$1 ( \2759 , \2758 , \1647 );
mnand \mul_18_12_g22320/U$1 ( \2760 , \2757 , \2759 );
mnand \mul_18_12_g23035/U$1 ( \2761 , \2753 , \2760 );
mnot \mul_18_12_g22258/U$2 ( \2762 , \2760 );
mnand \mul_18_12_g22258/U$1 ( \2763 , \2762 , \2752 );
mnand \mul_18_12_g22248/U$1 ( \2764 , \2761 , \2763 );
mnot \mul_18_12_g22232/U$3 ( \2765 , \2764 );
mand \mul_18_12_g2/U$1 ( \2766 , \1388 , \1657 , \1161 );
mnot \mul_18_12_g22234/U$3 ( \2767 , \2766 );
mnot \g37265/U$2 ( \2768 , \1530 );
mnot \mul_18_12_g22245/U$3 ( \2769 , \1539 );
mnand \mul_18_12_g22257/U$1 ( \2770 , \1309 , \1527 );
mnot \mul_18_12_g22245/U$4 ( \2771 , \2770 );
mor \mul_18_12_g22245/U$2 ( \2772 , \2769 , \2771 );
mnand \mul_18_12_g22245/U$1 ( \2773 , \2772 , \1214 );
mnand \g37265/U$1 ( \2774 , \2768 , \2773 );
mnot \mul_18_12_g22234/U$4 ( \2775 , \2774 );
mor \mul_18_12_g22234/U$2 ( \2776 , \2767 , \2775 );
mnot \mul_18_12_g22294/U$1 ( \2777 , \1543 );
mnot \g37117/U$3 ( \2778 , \2777 );
mnot \g37117/U$4 ( \2779 , \1657 );
mor \g37117/U$2 ( \2780 , \2778 , \2779 );
mnand \g37117/U$1 ( \2781 , \2780 , \1655 );
mnot \mul_18_12_g22259/U$1 ( \2782 , \2781 );
mnand \mul_18_12_g22234/U$1 ( \2783 , \2776 , \2782 );
mnot \mul_18_12_g22232/U$4 ( \2784 , \2783 );
mor \mul_18_12_g22232/U$2 ( \2785 , \2765 , \2784 );
mor \mul_18_12_g22232/U$5 ( \2786 , \2764 , \2783 );
mnand \mul_18_12_g22232/U$1 ( \2787 , \2785 , \2786 );
mnand \g4788/U$1 ( \2788 , \2787 , \1668 );
mnand \g4540/U$1 ( \2789 , \2475 , \a[14] );
mnand \g4516/U$1 ( \2790 , \2603 , \2657 , \2788 , \2789 );
mbuf \g4800/U$1 ( \2791 , \667 );
mor \g4784/U$1 ( \2792 , \a[11] , \b[11] );
mand \g4571/U$2 ( \2793 , \2791 , \2792 );
mand \g4786/U$1 ( \2794 , \b[11] , \c[11] );
mnot \g4586/U$3 ( \2795 , \2794 );
mnot \g4586/U$4 ( \2796 , \922 );
mor \g4586/U$2 ( \2797 , \2795 , \2796 );
mxor \g4731/U$1 ( \2798 , \c[11] , \d[11] );
mand \g4613/U$2 ( \2799 , \2615 , \2798 );
mnor \add_17_12_g6744/U$1 ( \2800 , \748 , \774 );
mnot \add_17_12_g6685/U$3 ( \2801 , \2800 );
mnot \add_17_12_g6779/U$1 ( \2802 , \749 );
mand \add_17_12_g6700/U$2 ( \2803 , \747 , \753 , \2802 );
mnot \add_17_12_g6721/U$3 ( \2804 , \2802 );
mnot \add_17_12_g6721/U$4 ( \2805 , \766 );
mor \add_17_12_g6721/U$2 ( \2806 , \2804 , \2805 );
mnand \add_17_12_g6721/U$1 ( \2807 , \2806 , \771 );
mnor \add_17_12_g6700/U$1 ( \2808 , \2803 , \2807 );
mnot \add_17_12_g6685/U$4 ( \2809 , \2808 );
mor \add_17_12_g6685/U$2 ( \2810 , \2801 , \2809 );
mor \add_17_12_g6685/U$5 ( \2811 , \2808 , \2800 );
mnand \add_17_12_g6685/U$1 ( \2812 , \2810 , \2811 );
mnot \g4626/U$3 ( \2813 , \2812 );
mnot \g4626/U$4 ( \2814 , \707 );
mor \g4626/U$2 ( \2815 , \2813 , \2814 );
mnor \add_16_12_g6744/U$1 ( \2816 , \833 , \859 );
mnot \add_16_12_g6685/U$3 ( \2817 , \2816 );
mnot \add_16_12_g6779/U$1 ( \2818 , \834 );
mand \add_16_12_g6700/U$2 ( \2819 , \832 , \838 , \2818 );
mnot \add_16_12_g6721/U$3 ( \2820 , \2818 );
mnot \add_16_12_g6721/U$4 ( \2821 , \851 );
mor \add_16_12_g6721/U$2 ( \2822 , \2820 , \2821 );
mnand \add_16_12_g6721/U$1 ( \2823 , \2822 , \856 );
mnor \add_16_12_g6700/U$1 ( \2824 , \2819 , \2823 );
mnot \add_16_12_g6685/U$4 ( \2825 , \2824 );
mor \add_16_12_g6685/U$2 ( \2826 , \2817 , \2825 );
mor \add_16_12_g6685/U$5 ( \2827 , \2824 , \2816 );
mnand \add_16_12_g6685/U$1 ( \2828 , \2826 , \2827 );
mand \g4649/U$2 ( \2829 , \880 , \2828 );
mnot \g4677/U$3 ( \2830 , \d[11] );
mnot \g4677/U$4 ( \2831 , \894 );
mor \g4677/U$2 ( \2832 , \2830 , \2831 );
mand \g4718/U$2 ( \2833 , \885 , \b[11] );
mand \g4718/U$3 ( \2834 , \909 , \c[11] );
mnor \g4718/U$1 ( \2835 , \2833 , \2834 );
mnand \g4677/U$1 ( \2836 , \2832 , \2835 );
mnor \g4649/U$1 ( \2837 , \2829 , \2836 );
mnand \g4626/U$1 ( \2838 , \2815 , \2837 );
mnor \g4613/U$1 ( \2839 , \2799 , \2838 );
mnand \g4586/U$1 ( \2840 , \2797 , \2839 );
mnor \g4571/U$1 ( \2841 , \2793 , \2840 );
mor \g36899/U$1 ( \2842 , \a[11] , \d[11] );
mbuf \g4837/U$1 ( \2843 , \648 );
mand \g36898/U$2 ( \2844 , \2842 , \2843 );
mnot \mul_18_12_g23038/U$2 ( \2845 , \1537 );
mnand \mul_18_12_g23038/U$1 ( \2846 , \2845 , \2770 );
mnot \mul_18_12_g22240/U$3 ( \2847 , \2846 );
mnot \mul_18_12_g22240/U$4 ( \2848 , \1214 );
mor \mul_18_12_g22240/U$2 ( \2849 , \2847 , \2848 );
mnot \mul_18_12_g22316/U$1 ( \2850 , \1538 );
mnand \mul_18_12_g22240/U$1 ( \2851 , \2849 , \2850 );
mnot \mul_18_12_g22272/U$2 ( \2852 , \1530 );
mnand \mul_18_12_g22272/U$1 ( \2853 , \2852 , \1541 );
mxor \g37039/U$1 ( \2854 , \2851 , \2853 );
mnor \g4735/U$1 ( \2855 , \2854 , \1667 );
mnor \g36898/U$1 ( \2856 , \2844 , \2855 );
mnand \g4902/U$1 ( \2857 , \2466 , \2474 );
mnot \g4562/U$1 ( \2858 , \2857 );
mbuf \g4561/U$1 ( \2859 , \2858 );
mnand \g4545/U$1 ( \2860 , \2859 , \a[11] );
mnot \mul_19_13_g22240/U$3 ( \2861 , \2285 );
mnot \mul_19_13_g23038/U$2 ( \2862 , \2280 );
mnand \mul_19_13_g23038/U$1 ( \2863 , \2862 , \2587 );
mnot \mul_19_13_g22240/U$4 ( \2864 , \2863 );
mor \mul_19_13_g22240/U$2 ( \2865 , \2861 , \2864 );
mnot \mul_19_13_g22316/U$1 ( \2866 , \2281 );
mnand \mul_19_13_g22240/U$1 ( \2867 , \2865 , \2866 );
mnot \mul_19_13_g22272/U$2 ( \2868 , \2273 );
mnand \mul_19_13_g22272/U$1 ( \2869 , \2868 , \2284 );
mnot \mul_19_13_g22271/U$1 ( \2870 , \2869 );
mand \mul_19_13_g22237/U$2 ( \2871 , \2867 , \2870 );
mnot \mul_19_13_g22237/U$4 ( \2872 , \2867 );
mand \mul_19_13_g22237/U$3 ( \2873 , \2872 , \2869 );
mnor \mul_19_13_g22237/U$1 ( \2874 , \2871 , \2873 );
mnand \g36905/U$1 ( \2875 , \2874 , \2413 );
mnand \g4517/U$1 ( \2876 , \2841 , \2856 , \2860 , \2875 );
mnot \g4799/U$1 ( \2877 , \666 );
mnot \g4656/U$3 ( \2878 , \2877 );
mnor \g4790/U$1 ( \2879 , \a[3] , \b[3] );
mnot \g4656/U$4 ( \2880 , \2879 );
mand \g4656/U$2 ( \2881 , \2878 , \2880 );
mnot \g4751/U$1 ( \2882 , \674 );
mand \g4656/U$5 ( \2883 , \648 , \2882 );
mnor \g4656/U$1 ( \2884 , \2881 , \2883 );
mnand \g4546/U$1 ( \2885 , \2858 , \a[3] );
mnot \g4863/U$1 ( \2886 , \921 );
mnot \g4862/U$1 ( \2887 , \2886 );
mand \g4755/U$1 ( \2888 , \b[3] , \c[3] );
mand \g4555/U$2 ( \2889 , \2887 , \2888 );
mxor \g4732/U$1 ( \2890 , \c[3] , \d[3] );
mnot \g4580/U$3 ( \2891 , \2890 );
mnot \g4580/U$4 ( \2892 , \697 );
mor \g4580/U$2 ( \2893 , \2891 , \2892 );
mnot \mul_19_13_g22437/U$3 ( \2894 , \2225 );
mnand \mul_19_13_g22493/U$1 ( \2895 , \2228 , \2204 );
mnot \mul_19_13_g22437/U$4 ( \2896 , \2895 );
mor \mul_19_13_g22437/U$2 ( \2897 , \2894 , \2896 );
mor \mul_19_13_g22437/U$5 ( \2898 , \2895 , \2225 );
mnand \mul_19_13_g22437/U$1 ( \2899 , \2897 , \2898 );
mand \g4596/U$2 ( \2900 , \2413 , \2899 );
mnot \mul_18_12_g22437/U$3 ( \2901 , \1507 );
mnand \mul_18_12_g22493/U$1 ( \2902 , \1487 , \1488 );
mnot \mul_18_12_g22437/U$4 ( \2903 , \2902 );
mor \mul_18_12_g22437/U$2 ( \2904 , \2901 , \2903 );
mor \mul_18_12_g22437/U$5 ( \2905 , \2902 , \1507 );
mnand \mul_18_12_g22437/U$1 ( \2906 , \2904 , \2905 );
mnot \g4609/U$3 ( \2907 , \2906 );
mnot \g4876/U$1 ( \2908 , \1667 );
mnot \g4609/U$4 ( \2909 , \2908 );
mor \g4609/U$2 ( \2910 , \2907 , \2909 );
mnot \add_17_12_g6757/U$2 ( \2911 , \732 );
mnand \add_17_12_g6757/U$1 ( \2912 , \2911 , \721 );
mnot \add_17_12_g6711/U$3 ( \2913 , \2912 );
mnand \add_17_12_g6717/U$1 ( \2914 , \720 , \722 );
mnot \add_17_12_g6711/U$4 ( \2915 , \2914 );
mor \add_17_12_g6711/U$2 ( \2916 , \2913 , \2915 );
mor \add_17_12_g6711/U$5 ( \2917 , \2914 , \2912 );
mnand \add_17_12_g6711/U$1 ( \2918 , \2916 , \2917 );
mand \g4627/U$2 ( \2919 , \707 , \2918 );
mnot \add_16_12_g6757/U$2 ( \2920 , \817 );
mnand \add_16_12_g6757/U$1 ( \2921 , \2920 , \806 );
mnot \add_16_12_g6711/U$3 ( \2922 , \2921 );
mnand \add_16_12_g6717/U$1 ( \2923 , \805 , \807 );
mnot \add_16_12_g6711/U$4 ( \2924 , \2923 );
mor \add_16_12_g6711/U$2 ( \2925 , \2922 , \2924 );
mor \add_16_12_g6711/U$5 ( \2926 , \2923 , \2921 );
mnand \add_16_12_g6711/U$1 ( \2927 , \2925 , \2926 );
mnot \g4634/U$3 ( \2928 , \2927 );
mnot \g4634/U$4 ( \2929 , \879 );
mor \g4634/U$2 ( \2930 , \2928 , \2929 );
mand \g4657/U$2 ( \2931 , \894 , \d[3] );
mnot \g4696/U$3 ( \2932 , \c[3] );
mnot \g4696/U$4 ( \2933 , \907 );
mor \g4696/U$2 ( \2934 , \2932 , \2933 );
mnand \g4747/U$1 ( \2935 , \885 , \b[3] );
mnand \g4696/U$1 ( \2936 , \2934 , \2935 );
mnor \g4657/U$1 ( \2937 , \2931 , \2936 );
mnand \g4634/U$1 ( \2938 , \2930 , \2937 );
mnor \g4627/U$1 ( \2939 , \2919 , \2938 );
mnand \g4609/U$1 ( \2940 , \2910 , \2939 );
mnor \g4596/U$1 ( \2941 , \2900 , \2940 );
mnand \g4580/U$1 ( \2942 , \2893 , \2941 );
mnor \g4555/U$1 ( \2943 , \2889 , \2942 );
mnand \g4519/U$1 ( \2944 , \2884 , \2885 , \2943 );
mbuf \g4518/U$1 ( \2945 , \2944 );
mnot \g4547/U$2 ( \2946 , \922 );
mand \g4558/U$1 ( \2947 , \2474 , \a[2] );
mnand \g4547/U$1 ( \2948 , \2946 , \2947 );
mand \g4738/U$1 ( \2949 , \b[2] , \c[2] );
mand \g4549/U$2 ( \2950 , \2887 , \2949 );
mxor \g4719/U$1 ( \2951 , \c[2] , \d[2] );
mnot \g4574/U$3 ( \2952 , \2951 );
mnot \g4574/U$4 ( \2953 , \2614 );
mor \g4574/U$2 ( \2954 , \2952 , \2953 );
mnot \mul_19_13_g22501/U$3 ( \2955 , \2222 );
mnot \mul_19_13_g22555/U$2 ( \2956 , \2224 );
mnor \mul_19_13_g22555/U$1 ( \2957 , \2956 , \2213 );
mnot \mul_19_13_g22501/U$4 ( \2958 , \2957 );
mor \mul_19_13_g22501/U$2 ( \2959 , \2955 , \2958 );
mor \mul_19_13_g22501/U$5 ( \2960 , \2957 , \2222 );
mnand \mul_19_13_g22501/U$1 ( \2961 , \2959 , \2960 );
mand \g4589/U$2 ( \2962 , \2413 , \2961 );
mnot \mul_18_12_g22501/U$3 ( \2963 , \1504 );
mnot \mul_18_12_g22555/U$2 ( \2964 , \1506 );
mnor \mul_18_12_g22555/U$1 ( \2965 , \2964 , \1496 );
mnot \mul_18_12_g22501/U$4 ( \2966 , \2965 );
mor \mul_18_12_g22501/U$2 ( \2967 , \2963 , \2966 );
mor \mul_18_12_g22501/U$5 ( \2968 , \2965 , \1504 );
mnand \mul_18_12_g22501/U$1 ( \2969 , \2967 , \2968 );
mnot \g4600/U$3 ( \2970 , \2969 );
mnot \g4600/U$4 ( \2971 , \2908 );
mor \g4600/U$2 ( \2972 , \2970 , \2971 );
mnand \add_17_12_g6748/U$1 ( \2973 , \719 , \722 );
mnot \add_17_12_g6716/U$3 ( \2974 , \2973 );
mnot \add_17_12_g6742/U$1 ( \2975 , \714 );
mnot \add_17_12_g6720/U$3 ( \2976 , \2975 );
mnot \add_17_12_g6720/U$4 ( \2977 , \717 );
mor \add_17_12_g6720/U$2 ( \2978 , \2976 , \2977 );
mnand \add_17_12_g6720/U$1 ( \2979 , \2978 , \715 );
mnot \add_17_12_g6716/U$4 ( \2980 , \2979 );
mor \add_17_12_g6716/U$2 ( \2981 , \2974 , \2980 );
mor \add_17_12_g6716/U$5 ( \2982 , \2979 , \2973 );
mnand \add_17_12_g6716/U$1 ( \2983 , \2981 , \2982 );
mand \g4614/U$2 ( \2984 , \707 , \2983 );
mnand \add_16_12_g6748/U$1 ( \2985 , \804 , \807 );
mnot \add_16_12_g6716/U$3 ( \2986 , \2985 );
mnot \add_16_12_g6742/U$1 ( \2987 , \799 );
mnot \add_16_12_g6720/U$3 ( \2988 , \2987 );
mnot \add_16_12_g6720/U$4 ( \2989 , \802 );
mor \add_16_12_g6720/U$2 ( \2990 , \2988 , \2989 );
mnand \add_16_12_g6720/U$1 ( \2991 , \2990 , \800 );
mnot \add_16_12_g6716/U$4 ( \2992 , \2991 );
mor \add_16_12_g6716/U$2 ( \2993 , \2986 , \2992 );
mor \add_16_12_g6716/U$5 ( \2994 , \2991 , \2985 );
mnand \add_16_12_g6716/U$1 ( \2995 , \2993 , \2994 );
mnot \g4635/U$3 ( \2996 , \2995 );
mnot \g4635/U$4 ( \2997 , \879 );
mor \g4635/U$2 ( \2998 , \2996 , \2997 );
mand \g4659/U$2 ( \2999 , \894 , \d[2] );
mnot \g4699/U$3 ( \3000 , \c[2] );
mnot \g4699/U$4 ( \3001 , \907 );
mor \g4699/U$2 ( \3002 , \3000 , \3001 );
mnand \g4746/U$1 ( \3003 , \885 , \b[2] );
mnand \g4699/U$1 ( \3004 , \3002 , \3003 );
mnor \g4659/U$1 ( \3005 , \2999 , \3004 );
mnand \g4635/U$1 ( \3006 , \2998 , \3005 );
mnor \g4614/U$1 ( \3007 , \2984 , \3006 );
mnand \g4600/U$1 ( \3008 , \2972 , \3007 );
mnor \g4589/U$1 ( \3009 , \2962 , \3008 );
mnand \g4574/U$1 ( \3010 , \2954 , \3009 );
mnor \g4549/U$1 ( \3011 , \2950 , \3010 );
mnot \g4910/U$2 ( \3012 , \683 );
mnand \g4910/U$1 ( \3013 , \3012 , \648 );
mor \g37051/U$2 ( \3014 , \b[2] , \a[2] );
mnand \g37051/U$1 ( \3015 , \3014 , \667 );
mnand \g4520/U$1 ( \3016 , \2948 , \3011 , \3013 , \3015 );
mand \g4741/U$1 ( \3017 , \b[1] , \c[1] );
mand \g4550/U$2 ( \3018 , \922 , \3017 );
mxor \g4721/U$1 ( \3019 , \c[1] , \d[1] );
mnot \g4575/U$3 ( \3020 , \3019 );
mnot \g4575/U$4 ( \3021 , \2614 );
mor \g4575/U$2 ( \3022 , \3020 , \3021 );
mor \mul_19_13_g23069/U$1 ( \3023 , \2219 , \2221 );
mand \mul_19_13_g22559/U$1 ( \3024 , \2222 , \3023 );
mand \g4590/U$2 ( \3025 , \2413 , \3024 );
mor \mul_18_12_g23069/U$1 ( \3026 , \1502 , \1503 );
mand \mul_18_12_g22559/U$1 ( \3027 , \1504 , \3026 );
mnot \g4601/U$3 ( \3028 , \3027 );
mnot \g4601/U$4 ( \3029 , \2908 );
mor \g4601/U$2 ( \3030 , \3028 , \3029 );
mnot \add_17_12_g6726/U$3 ( \3031 , \2975 );
mnand \add_17_12_g6762/U$1 ( \3032 , \717 , \715 );
mnot \add_17_12_g6726/U$4 ( \3033 , \3032 );
mor \add_17_12_g6726/U$2 ( \3034 , \3031 , \3033 );
mor \add_17_12_g6726/U$5 ( \3035 , \3032 , \2975 );
mnand \add_17_12_g6726/U$1 ( \3036 , \3034 , \3035 );
mand \g4617/U$2 ( \3037 , \707 , \3036 );
mnot \add_16_12_g6726/U$3 ( \3038 , \2987 );
mnand \add_16_12_g6762/U$1 ( \3039 , \802 , \800 );
mnot \add_16_12_g6726/U$4 ( \3040 , \3039 );
mor \add_16_12_g6726/U$2 ( \3041 , \3038 , \3040 );
mor \add_16_12_g6726/U$5 ( \3042 , \3039 , \2987 );
mnand \add_16_12_g6726/U$1 ( \3043 , \3041 , \3042 );
mnot \g4638/U$3 ( \3044 , \3043 );
mnot \g4638/U$4 ( \3045 , \879 );
mor \g4638/U$2 ( \3046 , \3044 , \3045 );
mand \g4658/U$2 ( \3047 , \894 , \d[1] );
mnot \g4701/U$3 ( \3048 , \c[1] );
mnot \g4701/U$4 ( \3049 , \907 );
mor \g4701/U$2 ( \3050 , \3048 , \3049 );
mnand \g4780/U$1 ( \3051 , \885 , \b[1] );
mnand \g4701/U$1 ( \3052 , \3050 , \3051 );
mnor \g4658/U$1 ( \3053 , \3047 , \3052 );
mnand \g4638/U$1 ( \3054 , \3046 , \3053 );
mnor \g4617/U$1 ( \3055 , \3037 , \3054 );
mnand \g4601/U$1 ( \3056 , \3030 , \3055 );
mnor \g4590/U$1 ( \3057 , \3025 , \3056 );
mnand \g4575/U$1 ( \3058 , \3022 , \3057 );
mnor \g4550/U$1 ( \3059 , \3018 , \3058 );
mand \g4559/U$1 ( \3060 , \2474 , \a[1] );
mnand \g4915/U$1 ( \3061 , \3060 , \2886 );
mnot \g4846/U$1 ( \3062 , \b[1] );
mnot \g4686/U$3 ( \3063 , \3062 );
mnot \g4817/U$1 ( \3064 , \a[1] );
mnot \g4686/U$4 ( \3065 , \3064 );
mor \g4686/U$2 ( \3066 , \3063 , \3065 );
mnand \g4686/U$1 ( \3067 , \3066 , \667 );
mnot \g4911/U$2 ( \3068 , \680 );
mnand \g4911/U$1 ( \3069 , \3068 , \648 );
mnand \g4521/U$1 ( \3070 , \3059 , \3061 , \3067 , \3069 );
mnot \g4522/U$3 ( \3071 , \a[8] );
mnot \g4566/U$1 ( \3072 , \2857 );
mnot \g36946/U$2 ( \3073 , \3072 );
mnor \g4793/U$1 ( \3074 , \648 , \666 );
mnand \g36946/U$1 ( \3075 , \3073 , \3074 );
mnot \g4522/U$4 ( \3076 , \3075 );
mor \g4522/U$2 ( \3077 , \3071 , \3076 );
mnot \g4688/U$3 ( \3078 , \c[8] );
mnot \g4688/U$4 ( \3079 , \922 );
mor \g4688/U$2 ( \3080 , \3078 , \3079 );
mnot \g4801/U$1 ( \3081 , \667 );
mnand \g4688/U$1 ( \3082 , \3080 , \3081 );
mand \g4557/U$2 ( \3083 , \3082 , \b[8] );
mnot \g4581/U$3 ( \3084 , \d[8] );
mnot \g4581/U$4 ( \3085 , \648 );
mor \g4581/U$2 ( \3086 , \3084 , \3085 );
mnot \mul_18_12_g22253/U$3 ( \3087 , \1527 );
mbuf \mul_18_12_g22336/U$1 ( \3088 , \1287 );
mbuf \mul_18_12_g22338/U$1 ( \3089 , \1534 );
mnand \mul_18_12_g23040/U$1 ( \3090 , \3088 , \3089 );
mnot \mul_18_12_g22253/U$4 ( \3091 , \3090 );
mor \mul_18_12_g22253/U$2 ( \3092 , \3087 , \3091 );
mor \mul_18_12_g22253/U$5 ( \3093 , \1528 , \3090 );
mnand \mul_18_12_g22253/U$1 ( \3094 , \3092 , \3093 );
mand \g4604/U$2 ( \3095 , \3094 , \2908 );
mnot \add_16_12_g6755/U$2 ( \3096 , \837 );
mnand \add_16_12_g6755/U$1 ( \3097 , \3096 , \848 );
mnot \add_16_12_g6701/U$3 ( \3098 , \3097 );
mnot \add_16_12_g6701/U$4 ( \3099 , \832 );
mor \add_16_12_g6701/U$2 ( \3100 , \3098 , \3099 );
mor \add_16_12_g6701/U$5 ( \3101 , \832 , \3097 );
mnand \add_16_12_g6701/U$1 ( \3102 , \3100 , \3101 );
mnot \g4642/U$3 ( \3103 , \3102 );
mnot \g4642/U$4 ( \3104 , \880 );
mor \g4642/U$2 ( \3105 , \3103 , \3104 );
mand \g37082/U$2 ( \3106 , \894 , \d[8] );
mand \g37082/U$3 ( \3107 , \c[8] , \909 );
mand \g37082/U$4 ( \3108 , \885 , \b[8] );
mnor \g37082/U$1 ( \3109 , \3106 , \3107 , \3108 );
mnand \g4642/U$1 ( \3110 , \3105 , \3109 );
mnot \g37215/U$2 ( \3111 , \3110 );
mnot \add_17_12_g6755/U$2 ( \3112 , \752 );
mnand \add_17_12_g6755/U$1 ( \3113 , \3112 , \763 );
mnot \add_17_12_g6701/U$3 ( \3114 , \3113 );
mnot \add_17_12_g6701/U$4 ( \3115 , \747 );
mor \add_17_12_g6701/U$2 ( \3116 , \3114 , \3115 );
mor \add_17_12_g6701/U$5 ( \3117 , \747 , \3113 );
mnand \add_17_12_g6701/U$1 ( \3118 , \3116 , \3117 );
mnand \g37216/U$1 ( \3119 , \3118 , \707 );
mnand \g37215/U$1 ( \3120 , \3111 , \3119 );
mnor \g4604/U$1 ( \3121 , \3095 , \3120 );
mxor \g4724/U$1 ( \3122 , \c[8] , \d[8] );
mnand \g4653/U$1 ( \3123 , \2614 , \3122 );
mbuf \mul_19_13_g22336/U$1 ( \3124 , \2027 );
mbuf \mul_19_13_g22338/U$1 ( \3125 , \2277 );
mnand \mul_19_13_g23040/U$1 ( \3126 , \3124 , \3125 );
mnot \mul_19_13_g22253/U$3 ( \3127 , \3126 );
mnot \mul_19_13_g22253/U$4 ( \3128 , \2270 );
mor \mul_19_13_g22253/U$2 ( \3129 , \3127 , \3128 );
mor \mul_19_13_g22253/U$5 ( \3130 , \2271 , \3126 );
mnand \mul_19_13_g22253/U$1 ( \3131 , \3129 , \3130 );
mnand \g4758/U$1 ( \3132 , \3131 , \2413 );
mand \g4583/U$1 ( \3133 , \3121 , \3123 , \3132 );
mnand \g4581/U$1 ( \3134 , \3086 , \3133 );
mnor \g4557/U$1 ( \3135 , \3083 , \3134 );
mnand \g4522/U$1 ( \3136 , \3077 , \3135 );
mnot \g4630/U$3 ( \3137 , \689 );
mnot \g4630/U$4 ( \3138 , \649 );
mor \g4630/U$2 ( \3139 , \3137 , \3138 );
mnot \g4671/U$3 ( \3140 , \b[12] );
mnot \g4671/U$4 ( \3141 , \922 );
mor \g4671/U$2 ( \3142 , \3140 , \3141 );
mand \g4693/U$2 ( \3143 , \697 , \687 );
mnor \g4693/U$1 ( \3144 , \3143 , \909 );
mnand \g4671/U$1 ( \3145 , \3142 , \3144 );
mnand \g4631/U$1 ( \3146 , \3145 , \c[12] );
mnand \g4630/U$1 ( \3147 , \3139 , \3146 );
mnand \g4544/U$1 ( \3148 , \2475 , \a[12] );
mnot \g4865/U$1 ( \3149 , \b[12] );
mnot \g4689/U$3 ( \3150 , \3149 );
mnot \g4689/U$4 ( \3151 , \688 );
mor \g4689/U$2 ( \3152 , \3150 , \3151 );
mnand \g4689/U$1 ( \3153 , \3152 , \667 );
mnot \g4857/U$1 ( \3154 , \c[12] );
mnot \g4694/U$3 ( \3155 , \3154 );
mnot \g4694/U$4 ( \3156 , \697 );
mor \g4694/U$2 ( \3157 , \3155 , \3156 );
mnand \g4694/U$1 ( \3158 , \3157 , \893 );
mand \g4632/U$2 ( \3159 , \3158 , \d[12] );
mnot \add_17_12_g6766/U$2 ( \3160 , \758 );
mnand \add_17_12_g6766/U$1 ( \3161 , \3160 , \779 );
mnot \add_17_12_g6690/U$3 ( \3162 , \3161 );
mnot \add_17_12_g6698/U$3 ( \3163 , \754 );
mnot \add_17_12_g6698/U$4 ( \3164 , \747 );
mor \add_17_12_g6698/U$2 ( \3165 , \3163 , \3164 );
mnand \add_17_12_g6698/U$1 ( \3166 , \3165 , \777 );
mnot \add_17_12_g6690/U$4 ( \3167 , \3166 );
mor \add_17_12_g6690/U$2 ( \3168 , \3162 , \3167 );
mor \add_17_12_g6690/U$5 ( \3169 , \3166 , \3161 );
mnand \add_17_12_g6690/U$1 ( \3170 , \3168 , \3169 );
mnot \g4673/U$3 ( \3171 , \3170 );
mnot \g4673/U$4 ( \3172 , \707 );
mor \g4673/U$2 ( \3173 , \3171 , \3172 );
mnot \g4714/U$3 ( \3174 , \886 );
mnot \g4714/U$4 ( \3175 , \3149 );
mand \g4714/U$2 ( \3176 , \3174 , \3175 );
mnot \add_16_12_g6766/U$2 ( \3177 , \843 );
mnand \add_16_12_g6766/U$1 ( \3178 , \3177 , \864 );
mnot \add_16_12_g6690/U$3 ( \3179 , \3178 );
mnot \add_16_12_g6698/U$3 ( \3180 , \839 );
mnot \add_16_12_g6698/U$4 ( \3181 , \832 );
mor \add_16_12_g6698/U$2 ( \3182 , \3180 , \3181 );
mnand \add_16_12_g6698/U$1 ( \3183 , \3182 , \862 );
mnot \add_16_12_g6690/U$4 ( \3184 , \3183 );
mor \add_16_12_g6690/U$2 ( \3185 , \3179 , \3184 );
mor \add_16_12_g6690/U$5 ( \3186 , \3183 , \3178 );
mnand \add_16_12_g6690/U$1 ( \3187 , \3185 , \3186 );
mand \g4714/U$5 ( \3188 , \880 , \3187 );
mnor \g4714/U$1 ( \3189 , \3176 , \3188 );
mnand \g4673/U$1 ( \3190 , \3173 , \3189 );
mnor \g4632/U$1 ( \3191 , \3159 , \3190 );
mnand \g4539/U$1 ( \3192 , \3148 , \3153 , \3191 );
mnor \g4524/U$1 ( \3193 , \3147 , \3192 );
mnot \g4525/U$3 ( \3194 , \a[0] );
mnot \g4556_dup/U$2 ( \3195 , \3072 );
mnand \g4556_dup/U$1 ( \3196 , \3195 , \3074 );
mnot \g4525/U$4 ( \3197 , \3196 );
mor \g4525/U$2 ( \3198 , \3194 , \3197 );
mnot \g4587/U$3 ( \3199 , \c[0] );
mnot \g4663/U$3 ( \3200 , \b[0] );
mnot \g4663/U$4 ( \3201 , \2887 );
mor \g4663/U$2 ( \3202 , \3200 , \3201 );
mnot \g4864/U$1 ( \3203 , \d[0] );
mand \g4695/U$2 ( \3204 , \903 , \3203 );
mnor \g4695/U$1 ( \3205 , \3204 , \909 );
mnand \g4663/U$1 ( \3206 , \3202 , \3205 );
mnot \g4587/U$4 ( \3207 , \3206 );
mor \g4587/U$2 ( \3208 , \3199 , \3207 );
mnot \g4856/U$1 ( \3209 , \c[0] );
mnot \g4691/U$3 ( \3210 , \3209 );
mnot \g4691/U$4 ( \3211 , \903 );
mor \g4691/U$2 ( \3212 , \3210 , \3211 );
mnand \g4691/U$1 ( \3213 , \3212 , \893 );
mand \g4598/U$2 ( \3214 , \3213 , \d[0] );
mnot \mul_19_13_g22976/U$1 ( \3215 , \2220 );
mnot \g4618/U$3 ( \3216 , \3215 );
mnot \g4618/U$4 ( \3217 , \2413 );
mor \g4618/U$2 ( \3218 , \3216 , \3217 );
mnot \mul_18_12_g22976/U$1 ( \3219 , \684 );
mand \g4639/U$2 ( \3220 , \1668 , \3219 );
mxor \add_17_12_g6768/U$1 ( \3221 , \b[0] , \d[0] );
mnot \g4664/U$3 ( \3222 , \3221 );
mnot \g4664/U$4 ( \3223 , \707 );
mor \g4664/U$2 ( \3224 , \3222 , \3223 );
mxor \add_16_12_g6768/U$1 ( \3225 , \a[0] , \c[0] );
mand \g4698/U$2 ( \3226 , \880 , \3225 );
mand \g4698/U$3 ( \3227 , \885 , \b[0] );
mnor \g4698/U$1 ( \3228 , \3226 , \3227 );
mnand \g4664/U$1 ( \3229 , \3224 , \3228 );
mnor \g4639/U$1 ( \3230 , \3220 , \3229 );
mnand \g4618/U$1 ( \3231 , \3218 , \3230 );
mnor \g4598/U$1 ( \3232 , \3214 , \3231 );
mnand \g4587/U$1 ( \3233 , \3208 , \3232 );
mnot \g4702/U$3 ( \3234 , \d[0] );
mbuf \g4838/U$1 ( \3235 , \648 );
mnot \g4702/U$4 ( \3236 , \3235 );
mor \g4702/U$2 ( \3237 , \3234 , \3236 );
mnand \g4778/U$1 ( \3238 , \2791 , \b[0] );
mnand \g4702/U$1 ( \3239 , \3237 , \3238 );
mnor \g4572/U$1 ( \3240 , \3233 , \3239 );
mnand \g4525/U$1 ( \3241 , \3198 , \3240 );
mnot \g4526/U$3 ( \3242 , \a[7] );
mnot \g4526/U$4 ( \3243 , \3075 );
mor \g4526/U$2 ( \3244 , \3242 , \3243 );
mnot \g4706/U$3 ( \3245 , \d[7] );
mnot \g4706/U$4 ( \3246 , \648 );
mor \g4706/U$2 ( \3247 , \3245 , \3246 );
mnand \g4768/U$1 ( \3248 , \667 , \b[7] );
mnand \g4706/U$1 ( \3249 , \3247 , \3248 );
mand \g4769/U$1 ( \3250 , \b[7] , \c[7] );
mnot \g4551/U$3 ( \3251 , \3250 );
mnot \g4551/U$4 ( \3252 , \922 );
mor \g4551/U$2 ( \3253 , \3251 , \3252 );
mxor \g4726/U$1 ( \3254 , \c[7] , \d[7] );
mand \g4576/U$2 ( \3255 , \2615 , \3254 );
mnand \mul_19_13_g23043/U$1 ( \3256 , \2269 , \2158 );
mxnor \g36566/U$1 ( \3257 , \2264 , \3256 );
mnot \g4592/U$3 ( \3258 , \3257 );
mnot \g4592/U$4 ( \3259 , \2413 );
mor \g4592/U$2 ( \3260 , \3258 , \3259 );
mbuf \mul_18_12_g22307/U$1 ( \3261 , \1523 );
mnot \mul_18_12_g22283/U$3 ( \3262 , \3261 );
mnand \mul_18_12_g23043/U$1 ( \3263 , \1526 , \1417 );
mnot \mul_18_12_g22283/U$4 ( \3264 , \3263 );
mor \mul_18_12_g22283/U$2 ( \3265 , \3262 , \3264 );
mor \mul_18_12_g22283/U$5 ( \3266 , \3263 , \3261 );
mnand \mul_18_12_g22283/U$1 ( \3267 , \3265 , \3266 );
mand \g4605/U$2 ( \3268 , \2908 , \3267 );
mnot \add_17_12_g2/U$2 ( \3269 , \729 );
mnand \add_17_12_g2/U$1 ( \3270 , \3269 , \736 );
mnot \add_17_12_g6691/U$3 ( \3271 , \3270 );
mnor \add_17_12_g6749/U$1 ( \3272 , \732 , \718 );
mand \add_17_12_g6713/U$2 ( \3273 , \2979 , \3272 );
mor \add_17_12_g6739/U$2 ( \3274 , \732 , \722 );
mnand \add_17_12_g6739/U$1 ( \3275 , \3274 , \721 );
mnor \add_17_12_g6713/U$1 ( \3276 , \3273 , \3275 );
mnot \add_17_12_g6730/U$2 ( \3277 , \728 );
mnand \add_17_12_g6730/U$1 ( \3278 , \3277 , \727 );
mor \add_17_12_g6704/U$2 ( \3279 , \3276 , \3278 );
mand \add_17_12_g6731/U$1 ( \3280 , \744 , \742 );
mor \add_17_12_g6704/U$3 ( \3281 , \728 , \3280 );
mnand \add_17_12_g6704/U$1 ( \3282 , \3279 , \3281 , \741 );
mnot \add_17_12_g6691/U$4 ( \3283 , \3282 );
mor \add_17_12_g6691/U$2 ( \3284 , \3271 , \3283 );
mor \add_17_12_g6691/U$5 ( \3285 , \3282 , \3270 );
mnand \add_17_12_g6691/U$1 ( \3286 , \3284 , \3285 );
mnot \g4622/U$3 ( \3287 , \3286 );
mnot \g4622/U$4 ( \3288 , \707 );
mor \g4622/U$2 ( \3289 , \3287 , \3288 );
mnot \add_16_12_g2/U$2 ( \3290 , \814 );
mnand \add_16_12_g2/U$1 ( \3291 , \3290 , \821 );
mnot \add_16_12_g6691/U$3 ( \3292 , \3291 );
mnor \add_16_12_g6749/U$1 ( \3293 , \817 , \803 );
mand \g37285/U$2 ( \3294 , \2991 , \3293 );
mor \add_16_12_g6739/U$2 ( \3295 , \817 , \807 );
mnand \add_16_12_g6739/U$1 ( \3296 , \3295 , \806 );
mnor \g37285/U$1 ( \3297 , \3294 , \3296 );
mnot \add_16_12_g6730/U$2 ( \3298 , \813 );
mnand \add_16_12_g6730/U$1 ( \3299 , \3298 , \812 );
mor \add_16_12_g6704/U$2 ( \3300 , \3297 , \3299 );
mand \add_16_12_g6731/U$1 ( \3301 , \829 , \827 );
mor \add_16_12_g6704/U$3 ( \3302 , \813 , \3301 );
mnand \add_16_12_g6704/U$1 ( \3303 , \3300 , \3302 , \826 );
mnot \add_16_12_g6691/U$4 ( \3304 , \3303 );
mor \add_16_12_g6691/U$2 ( \3305 , \3292 , \3304 );
mor \add_16_12_g6691/U$5 ( \3306 , \3303 , \3291 );
mnand \add_16_12_g6691/U$1 ( \3307 , \3305 , \3306 );
mand \g4645/U$2 ( \3308 , \880 , \3307 );
mnot \g4669/U$3 ( \3309 , \d[7] );
mnot \g4669/U$4 ( \3310 , \894 );
mor \g4669/U$2 ( \3311 , \3309 , \3310 );
mnot \g4709/U$3 ( \3312 , \886 );
mnot \g4844/U$1 ( \3313 , \b[7] );
mnot \g4709/U$4 ( \3314 , \3313 );
mand \g4709/U$2 ( \3315 , \3312 , \3314 );
mand \g4709/U$5 ( \3316 , \907 , \c[7] );
mnor \g4709/U$1 ( \3317 , \3315 , \3316 );
mnand \g4669/U$1 ( \3318 , \3311 , \3317 );
mnor \g4645/U$1 ( \3319 , \3308 , \3318 );
mnand \g4622/U$1 ( \3320 , \3289 , \3319 );
mnor \g4605/U$1 ( \3321 , \3268 , \3320 );
mnand \g4592/U$1 ( \3322 , \3260 , \3321 );
mnor \g4576/U$1 ( \3323 , \3255 , \3322 );
mnand \g4551/U$1 ( \3324 , \3253 , \3323 );
mnor \g4533/U$1 ( \3325 , \3249 , \3324 );
mnand \g4526/U$1 ( \3326 , \3244 , \3325 );
mnot \g4527/U$3 ( \3327 , \a[6] );
mnot \g4527/U$4 ( \3328 , \3196 );
mor \g4527/U$2 ( \3329 , \3327 , \3328 );
mnot \g4710/U$3 ( \3330 , \d[6] );
mnot \g4710/U$4 ( \3331 , \649 );
mor \g4710/U$2 ( \3332 , \3330 , \3331 );
mnand \g4748/U$1 ( \3333 , \667 , \b[6] );
mnand \g4710/U$1 ( \3334 , \3332 , \3333 );
mand \g4773/U$1 ( \3335 , \b[6] , \c[6] );
mnot \g4552/U$3 ( \3336 , \3335 );
mnot \g4552/U$4 ( \3337 , \922 );
mor \g4552/U$2 ( \3338 , \3336 , \3337 );
mxor \g4727/U$1 ( \3339 , \c[6] , \d[6] );
mand \g4577/U$2 ( \3340 , \903 , \3339 );
mxor \mul_19_13_g22308/U$1 ( \3341 , \2178 , \2180 );
mxor \mul_19_13_g22308/U$1_r1 ( \3342 , \3341 , \2261 );
mnot \g4593/U$3 ( \3343 , \3342 );
mnot \g4593/U$4 ( \3344 , \2413 );
mor \g4593/U$2 ( \3345 , \3343 , \3344 );
mxor \mul_18_12_g22308/U$1 ( \3346 , \1440 , \1442 );
mxor \mul_18_12_g22308/U$1_r1 ( \3347 , \3346 , \1520 );
mand \g4606/U$2 ( \3348 , \2908 , \3347 );
mnot \add_17_12_g6746/U$2 ( \3349 , \728 );
mnand \add_17_12_g6746/U$1 ( \3350 , \3349 , \741 );
mnot \add_17_12_g6692/U$3 ( \3351 , \3350 );
mnot \add_17_12_g6760/U$1 ( \3352 , \727 );
mor \add_17_12_g6705/U$2 ( \3353 , \3276 , \3352 );
mnand \add_17_12_g6705/U$1 ( \3354 , \3353 , \3280 );
mnot \add_17_12_g6692/U$4 ( \3355 , \3354 );
mor \add_17_12_g6692/U$2 ( \3356 , \3351 , \3355 );
mor \add_17_12_g6692/U$5 ( \3357 , \3354 , \3350 );
mnand \add_17_12_g6692/U$1 ( \3358 , \3356 , \3357 );
mnot \g4623/U$3 ( \3359 , \3358 );
mnot \g4623/U$4 ( \3360 , \707 );
mor \g4623/U$2 ( \3361 , \3359 , \3360 );
mnot \add_16_12_g6746/U$2 ( \3362 , \813 );
mnand \add_16_12_g6746/U$1 ( \3363 , \3362 , \826 );
mnot \add_16_12_g6692/U$3 ( \3364 , \3363 );
mnot \add_16_12_g6760/U$1 ( \3365 , \812 );
mor \add_16_12_g6705/U$2 ( \3366 , \3297 , \3365 );
mnand \add_16_12_g6705/U$1 ( \3367 , \3366 , \3301 );
mnot \add_16_12_g6692/U$4 ( \3368 , \3367 );
mor \add_16_12_g6692/U$2 ( \3369 , \3364 , \3368 );
mor \add_16_12_g6692/U$5 ( \3370 , \3367 , \3363 );
mnand \add_16_12_g6692/U$1 ( \3371 , \3369 , \3370 );
mand \g4646/U$2 ( \3372 , \880 , \3371 );
mnot \g4672/U$3 ( \3373 , \d[6] );
mnot \g4672/U$4 ( \3374 , \894 );
mor \g4672/U$2 ( \3375 , \3373 , \3374 );
mand \g4712/U$2 ( \3376 , \885 , \b[6] );
mand \g4712/U$3 ( \3377 , \909 , \c[6] );
mnor \g4712/U$1 ( \3378 , \3376 , \3377 );
mnand \g4672/U$1 ( \3379 , \3375 , \3378 );
mnor \g4646/U$1 ( \3380 , \3372 , \3379 );
mnand \g4623/U$1 ( \3381 , \3361 , \3380 );
mnor \g4606/U$1 ( \3382 , \3348 , \3381 );
mnand \g4593/U$1 ( \3383 , \3345 , \3382 );
mnor \g4577/U$1 ( \3384 , \3340 , \3383 );
mnand \g4552/U$1 ( \3385 , \3338 , \3384 );
mnor \g4534/U$1 ( \3386 , \3334 , \3385 );
mnand \g4527/U$1 ( \3387 , \3329 , \3386 );
mnot \g4528/U$3 ( \3388 , \a[5] );
mnot \g4528/U$4 ( \3389 , \3075 );
mor \g4528/U$2 ( \3390 , \3388 , \3389 );
mnot \g4713/U$3 ( \3391 , \d[5] );
mnot \g4713/U$4 ( \3392 , \649 );
mor \g4713/U$2 ( \3393 , \3391 , \3392 );
mnand \g4903/U$1 ( \3394 , \667 , \b[5] );
mnand \g4713/U$1 ( \3395 , \3393 , \3394 );
mand \g4767/U$1 ( \3396 , \b[5] , \c[5] );
mnot \g4553/U$3 ( \3397 , \3396 );
mnot \g4553/U$4 ( \3398 , \922 );
mor \g4553/U$2 ( \3399 , \3397 , \3398 );
mxor \g4728/U$1 ( \3400 , \c[5] , \d[5] );
mand \g4578/U$2 ( \3401 , \3400 , \903 );
mnot \mul_19_13_g22377/U$2 ( \3402 , \2258 );
mnand \mul_19_13_g22377/U$1 ( \3403 , \3402 , \2260 );
mxor \g36567/U$1 ( \3404 , \3403 , \2248 );
mnot \g4594/U$3 ( \3405 , \3404 );
mnot \g4594/U$4 ( \3406 , \2413 );
mor \g4594/U$2 ( \3407 , \3405 , \3406 );
mnot \mul_18_12_g22377/U$2 ( \3408 , \1466 );
mnand \mul_18_12_g22377/U$1 ( \3409 , \3408 , \1519 );
mxor \g37069/U$1 ( \3410 , \1517 , \3409 );
mand \g4607/U$2 ( \3411 , \2908 , \3410 );
mnot \add_17_12_g6754/U$2 ( \3412 , \725 );
mnand \add_17_12_g6754/U$1 ( \3413 , \3412 , \742 );
mnot \add_17_12_g6693/U$3 ( \3414 , \3413 );
mor \add_17_12_g6702/U$2 ( \3415 , \3276 , \726 );
mnand \add_17_12_g6702/U$1 ( \3416 , \3415 , \743 );
mnot \add_17_12_g6693/U$4 ( \3417 , \3416 );
mor \add_17_12_g6693/U$2 ( \3418 , \3414 , \3417 );
mor \add_17_12_g6693/U$5 ( \3419 , \3416 , \3413 );
mnand \add_17_12_g6693/U$1 ( \3420 , \3418 , \3419 );
mnot \g4624/U$3 ( \3421 , \3420 );
mnot \g4624/U$4 ( \3422 , \707 );
mor \g4624/U$2 ( \3423 , \3421 , \3422 );
mnot \add_16_12_g6754/U$2 ( \3424 , \810 );
mnand \add_16_12_g6754/U$1 ( \3425 , \3424 , \827 );
mnot \add_16_12_g6693/U$3 ( \3426 , \3425 );
mor \add_16_12_g6702/U$2 ( \3427 , \811 , \3297 );
mnand \add_16_12_g6702/U$1 ( \3428 , \3427 , \828 );
mnot \add_16_12_g6693/U$4 ( \3429 , \3428 );
mor \add_16_12_g6693/U$2 ( \3430 , \3426 , \3429 );
mor \add_16_12_g6693/U$5 ( \3431 , \3428 , \3425 );
mnand \add_16_12_g6693/U$1 ( \3432 , \3430 , \3431 );
mand \g4647/U$2 ( \3433 , \880 , \3432 );
mnot \g4674/U$3 ( \3434 , \d[5] );
mnot \g4674/U$4 ( \3435 , \894 );
mor \g4674/U$2 ( \3436 , \3434 , \3435 );
mand \g4715/U$2 ( \3437 , \885 , \b[5] );
mand \g4715/U$3 ( \3438 , \909 , \c[5] );
mnor \g4715/U$1 ( \3439 , \3437 , \3438 );
mnand \g4674/U$1 ( \3440 , \3436 , \3439 );
mnor \g4647/U$1 ( \3441 , \3433 , \3440 );
mnand \g4624/U$1 ( \3442 , \3423 , \3441 );
mnor \g4607/U$1 ( \3443 , \3411 , \3442 );
mnand \g4594/U$1 ( \3444 , \3407 , \3443 );
mnor \g4578/U$1 ( \3445 , \3401 , \3444 );
mnand \g4553/U$1 ( \3446 , \3399 , \3445 );
mnor \g4535/U$1 ( \3447 , \3395 , \3446 );
mnand \g4528/U$1 ( \3448 , \3390 , \3447 );
mnot \g4529/U$3 ( \3449 , \a[4] );
mnot \g4529/U$4 ( \3450 , \3075 );
mor \g4529/U$2 ( \3451 , \3449 , \3450 );
mnot \g4716/U$3 ( \3452 , \d[4] );
mnot \g4716/U$4 ( \3453 , \648 );
mor \g4716/U$2 ( \3454 , \3452 , \3453 );
mnand \g4781/U$1 ( \3455 , \667 , \b[4] );
mnand \g4716/U$1 ( \3456 , \3454 , \3455 );
mand \g4783/U$1 ( \3457 , \b[4] , \c[4] );
mnot \g4554/U$3 ( \3458 , \3457 );
mnot \g4554/U$4 ( \3459 , \2887 );
mor \g4554/U$2 ( \3460 , \3458 , \3459 );
mxor \g4730/U$1 ( \3461 , \c[4] , \d[4] );
mand \g4579/U$2 ( \3462 , \903 , \3461 );
mnot \mul_19_13_g22382/U$3 ( \3463 , \2229 );
mnot \mul_19_13_g23050/U$2 ( \3464 , \2247 );
mnand \mul_19_13_g23050/U$1 ( \3465 , \3464 , \2245 );
mnot \mul_19_13_g22382/U$4 ( \3466 , \3465 );
mor \mul_19_13_g22382/U$2 ( \3467 , \3463 , \3466 );
mor \mul_19_13_g22382/U$5 ( \3468 , \3465 , \2229 );
mnand \mul_19_13_g22382/U$1 ( \3469 , \3467 , \3468 );
mnot \g4595/U$3 ( \3470 , \3469 );
mnot \g4595/U$4 ( \3471 , \2413 );
mor \g4595/U$2 ( \3472 , \3470 , \3471 );
mnot \mul_18_12_g22382/U$3 ( \3473 , \1509 );
mnot \mul_18_12_g23050/U$2 ( \3474 , \1516 );
mnand \mul_18_12_g23050/U$1 ( \3475 , \3474 , \1514 );
mnot \mul_18_12_g22382/U$4 ( \3476 , \3475 );
mor \mul_18_12_g22382/U$2 ( \3477 , \3473 , \3476 );
mor \mul_18_12_g22382/U$5 ( \3478 , \3475 , \1509 );
mnand \mul_18_12_g22382/U$1 ( \3479 , \3477 , \3478 );
mand \g4608/U$2 ( \3480 , \2908 , \3479 );
mnot \add_17_12_g6756/U$2 ( \3481 , \743 );
mnor \add_17_12_g6756/U$1 ( \3482 , \3481 , \726 );
mnot \add_17_12_g6706/U$3 ( \3483 , \3482 );
mnot \add_17_12_g6706/U$4 ( \3484 , \3276 );
mor \add_17_12_g6706/U$2 ( \3485 , \3483 , \3484 );
mor \add_17_12_g6706/U$5 ( \3486 , \3276 , \3482 );
mnand \add_17_12_g6706/U$1 ( \3487 , \3485 , \3486 );
mnot \g4625/U$3 ( \3488 , \3487 );
mnot \g4625/U$4 ( \3489 , \707 );
mor \g4625/U$2 ( \3490 , \3488 , \3489 );
mnot \add_16_12_g6756/U$2 ( \3491 , \828 );
mnor \add_16_12_g6756/U$1 ( \3492 , \3491 , \811 );
mnot \add_16_12_g6706/U$3 ( \3493 , \3492 );
mnot \add_16_12_g6706/U$4 ( \3494 , \3297 );
mor \add_16_12_g6706/U$2 ( \3495 , \3493 , \3494 );
mor \add_16_12_g6706/U$5 ( \3496 , \3297 , \3492 );
mnand \add_16_12_g6706/U$1 ( \3497 , \3495 , \3496 );
mand \g4648/U$2 ( \3498 , \880 , \3497 );
mnot \g4676/U$3 ( \3499 , \d[4] );
mnot \g4676/U$4 ( \3500 , \894 );
mor \g4676/U$2 ( \3501 , \3499 , \3500 );
mnot \g4717/U$3 ( \3502 , \886 );
mnot \g4880/U$1 ( \3503 , \b[4] );
mnot \g4717/U$4 ( \3504 , \3503 );
mand \g4717/U$2 ( \3505 , \3502 , \3504 );
mand \g4717/U$5 ( \3506 , \907 , \c[4] );
mnor \g4717/U$1 ( \3507 , \3505 , \3506 );
mnand \g4676/U$1 ( \3508 , \3501 , \3507 );
mnor \g4648/U$1 ( \3509 , \3498 , \3508 );
mnand \g4625/U$1 ( \3510 , \3490 , \3509 );
mnor \g4608/U$1 ( \3511 , \3480 , \3510 );
mnand \g4595/U$1 ( \3512 , \3472 , \3511 );
mnor \g4579/U$1 ( \3513 , \3462 , \3512 );
mnand \g4554/U$1 ( \3514 , \3460 , \3513 );
mnor \g4536/U$1 ( \3515 , \3456 , \3514 );
mnand \g4529/U$1 ( \3516 , \3451 , \3515 );
mnand \g4531/U$1 ( \3517 , \3196 , \a[15] );
mnot \mul_19_13_g22303/U$2 ( \3518 , \2281 );
mnand \mul_19_13_g22303/U$1 ( \3519 , \3518 , \1954 );
mxnor \g36563/U$1 ( \3520 , \2863 , \3519 );
mand \g4697/U$2 ( \3521 , \3520 , \2413 );
mnot \mul_18_12_g22303/U$2 ( \3522 , \1538 );
mnand \mul_18_12_g22303/U$1 ( \3523 , \3522 , \1214 );
mnot \mul_18_12_g22243/U$3 ( \3524 , \3523 );
mnot \mul_18_12_g22243/U$4 ( \3525 , \2846 );
mor \mul_18_12_g22243/U$2 ( \3526 , \3524 , \3525 );
mor \mul_18_12_g22243/U$5 ( \3527 , \2846 , \3523 );
mnand \mul_18_12_g22243/U$1 ( \3528 , \3526 , \3527 );
mand \g4697/U$3 ( \3529 , \3528 , \1668 );
mnor \g4697/U$1 ( \3530 , \3521 , \3529 );
mand \g4739/U$1 ( \3531 , \b[10] , \c[10] );
mnand \g4690/U$1 ( \3532 , \922 , \3531 );
mxor \g4720/U$1 ( \3533 , \c[10] , \d[10] );
mand \g4610/U$2 ( \3534 , \2615 , \3533 );
mnot \add_17_12_g6747/U$2 ( \3535 , \771 );
mnor \add_17_12_g6747/U$1 ( \3536 , \3535 , \749 );
mnot \add_17_12_g6686/U$3 ( \3537 , \3536 );
mand \add_17_12_g6694/U$2 ( \3538 , \747 , \753 );
mnor \add_17_12_g6694/U$1 ( \3539 , \3538 , \766 );
mnot \add_17_12_g6686/U$4 ( \3540 , \3539 );
mor \add_17_12_g6686/U$2 ( \3541 , \3537 , \3540 );
mor \add_17_12_g6686/U$5 ( \3542 , \3539 , \3536 );
mnand \add_17_12_g6686/U$1 ( \3543 , \3541 , \3542 );
mnot \g4615/U$3 ( \3544 , \3543 );
mnot \g4615/U$4 ( \3545 , \707 );
mor \g4615/U$2 ( \3546 , \3544 , \3545 );
mnot \add_16_12_g6747/U$2 ( \3547 , \856 );
mnor \add_16_12_g6747/U$1 ( \3548 , \3547 , \834 );
mnot \add_16_12_g6686/U$3 ( \3549 , \3548 );
mand \add_16_12_g6694/U$2 ( \3550 , \832 , \838 );
mnor \add_16_12_g6694/U$1 ( \3551 , \3550 , \851 );
mnot \add_16_12_g6686/U$4 ( \3552 , \3551 );
mor \add_16_12_g6686/U$2 ( \3553 , \3549 , \3552 );
mor \add_16_12_g6686/U$5 ( \3554 , \3551 , \3548 );
mnand \add_16_12_g6686/U$1 ( \3555 , \3553 , \3554 );
mand \g4636/U$2 ( \3556 , \880 , \3555 );
mnot \g4660/U$3 ( \3557 , \d[10] );
mnot \g4660/U$4 ( \3558 , \894 );
mor \g4660/U$2 ( \3559 , \3557 , \3558 );
mand \g4700/U$2 ( \3560 , \885 , \b[10] );
mand \g4700/U$3 ( \3561 , \907 , \c[10] );
mnor \g4700/U$1 ( \3562 , \3560 , \3561 );
mnand \g4660/U$1 ( \3563 , \3559 , \3562 );
mnor \g4636/U$1 ( \3564 , \3556 , \3563 );
mnand \g4615/U$1 ( \3565 , \3546 , \3564 );
mnor \g4610/U$1 ( \3566 , \3534 , \3565 );
mand \g4570/U$1 ( \3567 , \3530 , \3532 , \3566 );
mnot \g2/U$2 ( \3568 , \672 );
mnand \g2/U$1 ( \3569 , \3568 , \3235 );
mnand \g4541/U$1 ( \3570 , \2859 , \a[10] );
mor \g4736/U$1 ( \3571 , \a[10] , \b[10] );
mnand \g4683/U$1 ( \3572 , \2791 , \3571 );
mnand \g4537/U$1 ( \3573 , \3567 , \3569 , \3570 , \3572 );
mand \g4787/U$1 ( \3574 , \b[9] , \c[9] );
mand \g4661/U$2 ( \3575 , \2887 , \3574 );
mnot \mul_19_13_g22251/U$3 ( \3576 , \3124 );
mnot \mul_19_13_g22251/U$4 ( \3577 , \2270 );
mor \mul_19_13_g22251/U$2 ( \3578 , \3576 , \3577 );
mnand \mul_19_13_g22251/U$1 ( \3579 , \3578 , \3125 );
mnot \mul_19_13_g22312/U$2 ( \3580 , \2048 );
mnand \mul_19_13_g22312/U$1 ( \3581 , \3580 , \2279 );
mxnor \g36564/U$1 ( \3582 , \3579 , \3581 );
mnot \g4913/U$2 ( \3583 , \3582 );
mnor \g4913/U$1 ( \3584 , \3583 , \2412 );
mnor \g4661/U$1 ( \3585 , \3575 , \3584 );
mor \g4766/U$1 ( \3586 , \a[9] , \b[9] );
mand \g4569/U$2 ( \3587 , \667 , \3586 );
mnot \mul_18_12_g22312/U$2 ( \3588 , \1308 );
mnand \mul_18_12_g22312/U$1 ( \3589 , \3588 , \1536 );
mnot \mul_18_12_g22244/U$3 ( \3590 , \3589 );
mnot \mul_18_12_g22251/U$3 ( \3591 , \3088 );
mnot \mul_18_12_g22251/U$4 ( \3592 , \1527 );
mor \mul_18_12_g22251/U$2 ( \3593 , \3591 , \3592 );
mnand \mul_18_12_g22251/U$1 ( \3594 , \3593 , \3089 );
mnot \mul_18_12_g22244/U$4 ( \3595 , \3594 );
mor \mul_18_12_g22244/U$2 ( \3596 , \3590 , \3595 );
mor \mul_18_12_g22244/U$5 ( \3597 , \3594 , \3589 );
mnand \mul_18_12_g22244/U$1 ( \3598 , \3596 , \3597 );
mnand \g4740/U$1 ( \3599 , \3598 , \1668 );
mxor \g4722/U$1 ( \3600 , \c[9] , \d[9] );
mnand \g4652/U$1 ( \3601 , \2614 , \3600 );
mnot \add_17_12_g6750/U$2 ( \3602 , \751 );
mnand \add_17_12_g6750/U$1 ( \3603 , \3602 , \765 );
mnot \add_17_12_g6687/U$3 ( \3604 , \3603 );
mnot \add_17_12_g6708/U$1 ( \3605 , \747 );
mor \add_17_12_g6697/U$2 ( \3606 , \3605 , \752 );
mnand \add_17_12_g6697/U$1 ( \3607 , \3606 , \763 );
mnot \add_17_12_g6687/U$4 ( \3608 , \3607 );
mor \add_17_12_g6687/U$2 ( \3609 , \3604 , \3608 );
mor \add_17_12_g6687/U$5 ( \3610 , \3607 , \3603 );
mnand \add_17_12_g6687/U$1 ( \3611 , \3609 , \3610 );
mand \g4619/U$2 ( \3612 , \707 , \3611 );
mnot \add_16_12_g6750/U$2 ( \3613 , \836 );
mnand \add_16_12_g6750/U$1 ( \3614 , \3613 , \850 );
mnot \add_16_12_g6687/U$3 ( \3615 , \3614 );
mnot \fopt36961/U$1 ( \3616 , \832 );
mor \add_16_12_g6697/U$2 ( \3617 , \3616 , \837 );
mnand \add_16_12_g6697/U$1 ( \3618 , \3617 , \848 );
mnot \add_16_12_g6687/U$4 ( \3619 , \3618 );
mor \add_16_12_g6687/U$2 ( \3620 , \3615 , \3619 );
mor \add_16_12_g6687/U$5 ( \3621 , \3618 , \3614 );
mnand \add_16_12_g6687/U$1 ( \3622 , \3620 , \3621 );
mnot \g4640/U$3 ( \3623 , \3622 );
mnot \g4640/U$4 ( \3624 , \880 );
mor \g4640/U$2 ( \3625 , \3623 , \3624 );
mand \g37268/U$2 ( \3626 , \894 , \d[9] );
mand \g37268/U$3 ( \3627 , \b[9] , \885 );
mand \g37268/U$4 ( \3628 , \907 , \c[9] );
mnor \g37268/U$1 ( \3629 , \3626 , \3627 , \3628 );
mnand \g4640/U$1 ( \3630 , \3625 , \3629 );
mnor \g4619/U$1 ( \3631 , \3612 , \3630 );
mnand \g4591/U$1 ( \3632 , \3599 , \3601 , \3631 );
mnor \g4569/U$1 ( \3633 , \3587 , \3632 );
mnand \g4542/U$1 ( \3634 , \2858 , \a[9] );
mnot \g4762/U$1 ( \3635 , \673 );
mnand \g4682/U$1 ( \3636 , \2843 , \3635 );
mnand \g4538/U$1 ( \3637 , \3585 , \3633 , \3634 , \3636 );
mnot \mul_19_13_g22270/U$2 ( \3638 , \2129 );
mnor \mul_19_13_g22270/U$1 ( \3639 , \3638 , \2287 );
mnot \mul_19_13_g22233/U$3 ( \3640 , \3639 );
mnand \mul_19_13_g22238/U$1 ( \3641 , \2592 , \2284 );
mnot \mul_19_13_g22233/U$4 ( \3642 , \3641 );
mor \mul_19_13_g22233/U$2 ( \3643 , \3640 , \3642 );
mor \mul_19_13_g22233/U$5 ( \3644 , \3641 , \3639 );
mnand \mul_19_13_g22233/U$1 ( \3645 , \3643 , \3644 );
mand \g4708/U$2 ( \3646 , \3645 , \2413 );
mnot \mul_18_12_g22270/U$2 ( \3647 , \1388 );
mnor \mul_18_12_g22270/U$1 ( \3648 , \3647 , \2777 );
mnot \mul_18_12_g22233/U$3 ( \3649 , \3648 );
mnand \mul_18_12_g22238/U$1 ( \3650 , \2774 , \1541 );
mnot \mul_18_12_g22233/U$4 ( \3651 , \3650 );
mor \mul_18_12_g22233/U$2 ( \3652 , \3649 , \3651 );
mor \mul_18_12_g22233/U$5 ( \3653 , \3650 , \3648 );
mnand \mul_18_12_g22233/U$1 ( \3654 , \3652 , \3653 );
mand \g4708/U$3 ( \3655 , \3654 , \1668 );
mnor \g4708/U$1 ( \3656 , \3646 , \3655 );
mand \mul_18_12_g22246/U$1 ( \3657 , \2763 , \1657 , \1541 );
mand \mul_18_12_g22250/U$1 ( \3658 , \1539 , \2770 );
mnand \mul_18_12_g22276/U$1 ( \3659 , \1388 , \1214 );
mor \mul_18_12_g22239/U$2 ( \3660 , \3658 , \3659 );
mnand \mul_18_12_g22275/U$1 ( \3661 , \1388 , \1530 );
mnand \mul_18_12_g22239/U$1 ( \3662 , \3660 , \3661 );
mand \mul_18_12_g22235/U$2 ( \3663 , \3657 , \3662 );
mnot \mul_18_12_g22247/U$3 ( \3664 , \2781 );
mnot \mul_18_12_g22247/U$4 ( \3665 , \2763 );
mor \mul_18_12_g22247/U$2 ( \3666 , \3664 , \3665 );
mnand \mul_18_12_g22247/U$1 ( \3667 , \3666 , \2761 );
mnor \mul_18_12_g22235/U$1 ( \3668 , \3663 , \3667 );
mnot \fopt36737/U$1 ( \3669 , \2737 );
mnot \mul_18_12_g22298/U$3 ( \3670 , \3669 );
mnot \mul_18_12_g22298/U$4 ( \3671 , \2709 );
mor \mul_18_12_g22298/U$2 ( \3672 , \3670 , \3671 );
mnand \mul_18_12_g22298/U$1 ( \3673 , \3672 , \2748 );
mnot \mul_18_12_g23039/U$2 ( \3674 , \2709 );
mnand \mul_18_12_g23039/U$1 ( \3675 , \3674 , \2737 );
mnand \mul_18_12_g22282/U$1 ( \3676 , \3673 , \3675 );
mnot \g36897/U$3 ( \3677 , \2708 );
mnand \mul_18_12_g22403/U$1 ( \3678 , \2674 , \2697 );
mnot \g36897/U$4 ( \3679 , \3678 );
mor \g36897/U$2 ( \3680 , \3677 , \3679 );
mnot \mul_18_12_g23047/U$2 ( \3681 , \2674 );
mnand \mul_18_12_g23047/U$1 ( \3682 , \3681 , \2696 );
mnand \g36897/U$1 ( \3683 , \3680 , \3682 );
mnot \mul_18_12_g22654/U$3 ( \3684 , \2693 );
mnot \mul_18_12_g22654/U$4 ( \3685 , \1312 );
mor \mul_18_12_g22654/U$2 ( \3686 , \3684 , \3685 );
mxor \mul_18_12_g23080/U$1 ( \3687 , \d[5] , \a[11] );
mnand \mul_18_12_g22715/U$1 ( \3688 , \936 , \3687 );
mnand \mul_18_12_g22654/U$1 ( \3689 , \3686 , \3688 );
mand \g37126/U$2 ( \3690 , \1366 , \2671 );
mxor \g36641/U$1 ( \3691 , \d[11] , \a[5] );
mand \g37126/U$3 ( \3692 , \947 , \3691 );
mnor \g37126/U$1 ( \3693 , \3690 , \3692 );
mxor \g37120/U$1 ( \3694 , \3689 , \3693 );
mnot \mul_18_12_g22436/U$3 ( \3695 , \2664 );
mnot \mul_18_12_g22539/U$1 ( \3696 , \2666 );
mnot \mul_18_12_g22436/U$4 ( \3697 , \3696 );
mor \mul_18_12_g22436/U$2 ( \3698 , \3695 , \3697 );
mnot \mul_18_12_g22607/U$1 ( \3699 , \2664 );
mnot \mul_18_12_g22450/U$3 ( \3700 , \3699 );
mnot \mul_18_12_g22450/U$4 ( \3701 , \2666 );
mor \mul_18_12_g22450/U$2 ( \3702 , \3700 , \3701 );
mnand \mul_18_12_g22450/U$1 ( \3703 , \3702 , \2673 );
mnand \mul_18_12_g22436/U$1 ( \3704 , \3698 , \3703 );
mxnor \g37120/U$1_r1 ( \3705 , \3694 , \3704 );
mxor \mul_18_12_g22485/U$4 ( \3706 , \2716 , \2722 );
mand \mul_18_12_g22485/U$3 ( \3707 , \3706 , \2729 );
mand \mul_18_12_g22485/U$5 ( \3708 , \2716 , \2722 );
mor \mul_18_12_g22485/U$2 ( \3709 , \3707 , \3708 );
mand \mul_18_12_g22610/U$2 ( \3710 , \1583 , \2662 );
mxor \g36644/U$1 ( \3711 , \d[13] , \a[3] );
mand \mul_18_12_g22610/U$3 ( \3712 , \1335 , \3711 );
mnor \mul_18_12_g22610/U$1 ( \3713 , \3710 , \3712 );
mxor \mul_18_12_g22918/U$1 ( \3714 , \d[15] , \d[14] );
mxor \mul_18_12_g22874/U$1 ( \3715 , \a[0] , \d[15] );
mnand \mul_18_12_g22769/U$1 ( \3716 , \3714 , \3715 );
mor \mul_18_12_g22596/U$2 ( \3717 , \3716 , \2715 );
mxor \mul_18_12_g22889/U$1 ( \3718 , \a[1] , \d[15] );
mnand \mul_18_12_g22709/U$1 ( \3719 , \2715 , \3718 );
mnand \mul_18_12_g22596/U$1 ( \3720 , \3717 , \3719 );
mxor \g37130/U$1 ( \3721 , \3713 , \3720 );
mnot \mul_18_12_g22636/U$3 ( \3722 , \2686 );
mnot \mul_18_12_g22636/U$4 ( \3723 , \999 );
mor \mul_18_12_g22636/U$2 ( \3724 , \3722 , \3723 );
mnot \mul_18_12_g22962/U$2 ( \3725 , \d[7] );
mnand \mul_18_12_g22962/U$1 ( \3726 , \3725 , \a[9] );
mnot \mul_18_12_g22714/U$3 ( \3727 , \3726 );
mnot \mul_18_12_g23078/U$2 ( \3728 , \a[9] );
mnand \mul_18_12_g23078/U$1 ( \3729 , \3728 , \d[7] );
mnot \mul_18_12_g22714/U$4 ( \3730 , \3729 );
mor \mul_18_12_g22714/U$2 ( \3731 , \3727 , \3730 );
mnand \mul_18_12_g22714/U$1 ( \3732 , \3731 , \1003 );
mnand \mul_18_12_g22636/U$1 ( \3733 , \3724 , \3732 );
mxnor \g37130/U$1_r1 ( \3734 , \3721 , \3733 );
mnot \mul_18_12_g37186/U$2 ( \3735 , \3734 );
mxor \mul_18_12_g37186/U$1 ( \3736 , \3709 , \3735 );
mxor \mul_18_12_g23049/U$1 ( \3737 , \3705 , \3736 );
mxor \g36896/U$1 ( \3738 , \3683 , \3737 );
mnot \mul_18_12_g22574/U$3 ( \3739 , \2680 );
mnot \mul_18_12_g22574/U$4 ( \3740 , \1026 );
mor \mul_18_12_g22574/U$2 ( \3741 , \3739 , \3740 );
mxor \mul_18_12_g22906/U$1 ( \3742 , \d[9] , \a[7] );
mnand \mul_18_12_g22671/U$1 ( \3743 , \1058 , \3742 );
mnand \mul_18_12_g22574/U$1 ( \3744 , \3741 , \3743 );
mnot \mul_18_12_g22668/U$3 ( \3745 , \2727 );
mnot \mul_18_12_g22668/U$4 ( \3746 , \962 );
mor \mul_18_12_g22668/U$2 ( \3747 , \3745 , \3746 );
mxor \mul_18_12_g23079/U$1 ( \3748 , \d[3] , \a[13] );
mnand \mul_18_12_g22790/U$1 ( \3749 , \965 , \3748 );
mnand \mul_18_12_g22668/U$1 ( \3750 , \3747 , \3749 );
mxor \mul_18_12_g23066/U$1 ( \3751 , \3744 , \3750 );
mand \mul_18_12_g22702/U$2 ( \3752 , \1065 , \2720 );
mnot \mul_18_12_g22781/U$2 ( \3753 , \d[0] );
mxnor \mul_18_12_g23077/U$1 ( \3754 , \d[1] , \a[15] );
mnor \mul_18_12_g22781/U$1 ( \3755 , \3753 , \3754 );
mnor \mul_18_12_g22702/U$1 ( \3756 , \3752 , \3755 );
mnot \mul_18_12_g22575/U$3 ( \3757 , \3756 );
mor \mul_18_12_g22816/U$2 ( \3758 , \a[0] , \d[14] );
mnand \mul_18_12_g22816/U$1 ( \3759 , \3758 , \d[13] );
mnand \mul_18_12_g22952/U$1 ( \3760 , \a[0] , \d[14] );
mand \mul_18_12_g22806/U$1 ( \3761 , \3759 , \3760 , \d[15] );
mnot \mul_18_12_g22575/U$4 ( \3762 , \3761 );
mand \mul_18_12_g22575/U$2 ( \3763 , \3757 , \3762 );
mand \mul_18_12_g22575/U$5 ( \3764 , \3756 , \3761 );
mnor \mul_18_12_g22575/U$1 ( \3765 , \3763 , \3764 );
mxnor \mul_18_12_g23066/U$1_r1 ( \3766 , \3751 , \3765 );
mxor \mul_18_12_g22463/U$4 ( \3767 , \2682 , \2688 );
mand \mul_18_12_g22463/U$3 ( \3768 , \3767 , \2695 );
mand \mul_18_12_g22463/U$5 ( \3769 , \2682 , \2688 );
mor \mul_18_12_g22463/U$2 ( \3770 , \3768 , \3769 );
mxnor \mul_18_12_g23051/U$1 ( \3771 , \3766 , \3770 );
mnot \mul_18_12_g22345/U$3 ( \3772 , \3771 );
mxor \mul_18_12_g22369/U$4 ( \3773 , \2714 , \2730 );
mand \mul_18_12_g22369/U$3 ( \3774 , \3773 , \2736 );
mand \mul_18_12_g22369/U$5 ( \3775 , \2714 , \2730 );
mor \mul_18_12_g22369/U$2 ( \3776 , \3774 , \3775 );
mnot \mul_18_12_g22345/U$4 ( \3777 , \3776 );
mand \mul_18_12_g22345/U$2 ( \3778 , \3772 , \3777 );
mand \mul_18_12_g22345/U$5 ( \3779 , \3776 , \3771 );
mnor \mul_18_12_g22345/U$1 ( \3780 , \3778 , \3779 );
mxnor \g36896/U$1_r1 ( \3781 , \3738 , \3780 );
mxnor \mul_18_12_g23036/U$1 ( \3782 , \3676 , \3781 );
mnot \mul_18_12_g22254/U$1 ( \3783 , \3782 );
mand \mul_18_12_g22231/U$2 ( \3784 , \3668 , \3783 );
mnot \mul_18_12_g22231/U$4 ( \3785 , \3668 );
mand \mul_18_12_g22231/U$3 ( \3786 , \3785 , \3782 );
mnor \mul_18_12_g22231/U$1 ( \3787 , \3784 , \3786 );
mnand \g4749/U$1 ( \3788 , \3787 , \1668 );
mnot \g37196/U$2 ( \3789 , \2581 );
mnand \g37197/U$1 ( \3790 , \2403 , \2284 );
mnor \g37196/U$1 ( \3791 , \3789 , \3790 );
mand \mul_19_13_g22250/U$1 ( \3792 , \2282 , \2587 );
mnand \mul_19_13_g22276/U$1 ( \3793 , \2129 , \2285 );
mor \mul_19_13_g22239/U$2 ( \3794 , \3792 , \3793 );
mnand \mul_19_13_g22275/U$1 ( \3795 , \2129 , \2273 );
mnand \mul_19_13_g22239/U$1 ( \3796 , \3794 , \3795 );
mand \mul_19_13_g22235/U$2 ( \3797 , \3791 , \3796 );
mnot \mul_19_13_g22247/U$3 ( \3798 , \2596 );
mnot \mul_19_13_g22247/U$4 ( \3799 , \2581 );
mor \mul_19_13_g22247/U$2 ( \3800 , \3798 , \3799 );
mnand \mul_19_13_g22247/U$1 ( \3801 , \3800 , \2579 );
mnor \mul_19_13_g22235/U$1 ( \3802 , \3797 , \3801 );
mnot \mul_19_13_g22368/U$1 ( \3803 , \2555 );
mnot \mul_19_13_g22298/U$3 ( \3804 , \3803 );
mnot \mul_19_13_g22298/U$4 ( \3805 , \2528 );
mor \mul_19_13_g22298/U$2 ( \3806 , \3804 , \3805 );
mnand \mul_19_13_g22298/U$1 ( \3807 , \3806 , \2566 );
mnot \mul_19_13_g23039/U$2 ( \3808 , \2528 );
mnand \mul_19_13_g23039/U$1 ( \3809 , \3808 , \2555 );
mnand \mul_19_13_g22282/U$1 ( \3810 , \3807 , \3809 );
mnot \mul_19_13_g22574/U$3 ( \3811 , \2497 );
mnot \mul_19_13_g22574/U$4 ( \3812 , \1770 );
mor \mul_19_13_g22574/U$2 ( \3813 , \3811 , \3812 );
mxor \mul_19_13_g22906/U$1 ( \3814 , \c[9] , \b[7] );
mnand \mul_19_13_g22671/U$1 ( \3815 , \1802 , \3814 );
mnand \mul_19_13_g22574/U$1 ( \3816 , \3813 , \3815 );
mnot \mul_19_13_g22668/U$3 ( \3817 , \2546 );
mnot \mul_19_13_g22668/U$4 ( \3818 , \2370 );
mor \mul_19_13_g22668/U$2 ( \3819 , \3817 , \3818 );
mxor \mul_19_13_g23079/U$1 ( \3820 , \c[3] , \b[13] );
mnand \mul_19_13_g22790/U$1 ( \3821 , \1708 , \3820 );
mnand \mul_19_13_g22668/U$1 ( \3822 , \3819 , \3821 );
mxor \mul_19_13_g23066/U$1 ( \3823 , \3816 , \3822 );
mand \mul_19_13_g22702/U$2 ( \3824 , \1756 , \2539 );
mnot \mul_19_13_g22781/U$2 ( \3825 , \c[0] );
mxnor \mul_19_13_g23077/U$1 ( \3826 , \c[1] , \b[15] );
mnor \mul_19_13_g22781/U$1 ( \3827 , \3825 , \3826 );
mnor \mul_19_13_g22702/U$1 ( \3828 , \3824 , \3827 );
mnot \mul_19_13_g22575/U$3 ( \3829 , \3828 );
mor \mul_19_13_g22816/U$2 ( \3830 , \b[0] , \c[14] );
mnand \mul_19_13_g22816/U$1 ( \3831 , \3830 , \c[13] );
mnand \mul_19_13_g22952/U$1 ( \3832 , \b[0] , \c[14] );
mand \mul_19_13_g22806/U$1 ( \3833 , \3831 , \3832 , \c[15] );
mnot \mul_19_13_g22575/U$4 ( \3834 , \3833 );
mand \mul_19_13_g22575/U$2 ( \3835 , \3829 , \3834 );
mand \mul_19_13_g22575/U$5 ( \3836 , \3828 , \3833 );
mnor \mul_19_13_g22575/U$1 ( \3837 , \3835 , \3836 );
mxnor \mul_19_13_g23066/U$1_r1 ( \3838 , \3823 , \3837 );
mxor \mul_19_13_g22463/U$4 ( \3839 , \2501 , \2507 );
mand \mul_19_13_g22463/U$3 ( \3840 , \3839 , \2514 );
mand \mul_19_13_g22463/U$5 ( \3841 , \2501 , \2507 );
mor \mul_19_13_g22463/U$2 ( \3842 , \3840 , \3841 );
mxnor \mul_19_13_g23051/U$1 ( \3843 , \3838 , \3842 );
mnot \mul_19_13_g22345/U$3 ( \3844 , \3843 );
mxor \mul_19_13_g22369/U$4 ( \3845 , \2533 , \2549 );
mand \mul_19_13_g22369/U$3 ( \3846 , \3845 , \2554 );
mand \mul_19_13_g22369/U$5 ( \3847 , \2533 , \2549 );
mor \mul_19_13_g22369/U$2 ( \3848 , \3846 , \3847 );
mnot \mul_19_13_g22345/U$4 ( \3849 , \3848 );
mand \mul_19_13_g22345/U$2 ( \3850 , \3844 , \3849 );
mand \mul_19_13_g22345/U$5 ( \3851 , \3848 , \3843 );
mnor \mul_19_13_g22345/U$1 ( \3852 , \3850 , \3851 );
mnand \mul_19_13_g22403/U$1 ( \3853 , \2493 , \2516 );
mnot \mul_19_13_g22342/U$3 ( \3854 , \3853 );
mnot \mul_19_13_g22342/U$4 ( \3855 , \2527 );
mor \mul_19_13_g22342/U$2 ( \3856 , \3854 , \3855 );
mnot \mul_19_13_g23047/U$2 ( \3857 , \2493 );
mnand \mul_19_13_g23047/U$1 ( \3858 , \3857 , \2515 );
mnand \mul_19_13_g22342/U$1 ( \3859 , \3856 , \3858 );
mnot \mul_19_13_g22654/U$3 ( \3860 , \2512 );
mnot \mul_19_13_g22654/U$4 ( \3861 , \2052 );
mor \mul_19_13_g22654/U$2 ( \3862 , \3860 , \3861 );
mxor \mul_19_13_g23080/U$1 ( \3863 , \c[5] , \b[11] );
mnand \mul_19_13_g22715/U$1 ( \3864 , \1678 , \3863 );
mnand \mul_19_13_g22654/U$1 ( \3865 , \3862 , \3864 );
mnot \mul_19_13_g22548/U$3 ( \3866 , \3865 );
mand \g37109/U$2 ( \3867 , \2107 , \2490 );
mxor \g36602/U$1 ( \3868 , \c[11] , \b[5] );
mand \g37109/U$3 ( \3869 , \1689 , \3868 );
mnor \g37109/U$1 ( \3870 , \3867 , \3869 );
mnot \mul_19_13_g22548/U$4 ( \3871 , \3870 );
mand \mul_19_13_g22548/U$2 ( \3872 , \3866 , \3871 );
mand \mul_19_13_g22548/U$5 ( \3873 , \3865 , \3870 );
mnor \mul_19_13_g22548/U$1 ( \3874 , \3872 , \3873 );
mnot \mul_19_13_g22436/U$3 ( \3875 , \2483 );
mnot \mul_19_13_g22539/U$1 ( \3876 , \2485 );
mnot \mul_19_13_g22436/U$4 ( \3877 , \3876 );
mor \mul_19_13_g22436/U$2 ( \3878 , \3875 , \3877 );
mnot \mul_19_13_g22607/U$1 ( \3879 , \2483 );
mnot \mul_19_13_g22450/U$3 ( \3880 , \3879 );
mnot \mul_19_13_g22450/U$4 ( \3881 , \2485 );
mor \mul_19_13_g22450/U$2 ( \3882 , \3880 , \3881 );
mnand \mul_19_13_g22450/U$1 ( \3883 , \3882 , \2492 );
mnand \mul_19_13_g22436/U$1 ( \3884 , \3878 , \3883 );
mxor \g37113/U$1 ( \3885 , \3874 , \3884 );
mxor \mul_19_13_g22485/U$4 ( \3886 , \2535 , \2541 );
mand \mul_19_13_g22485/U$3 ( \3887 , \3886 , \2548 );
mand \mul_19_13_g22485/U$5 ( \3888 , \2535 , \2541 );
mor \mul_19_13_g22485/U$2 ( \3889 , \3887 , \3888 );
mand \mul_19_13_g22610/U$2 ( \3890 , \2341 , \2481 );
mxor \g36605/U$1 ( \3891 , \c[13] , \b[3] );
mand \mul_19_13_g22610/U$3 ( \3892 , \2075 , \3891 );
mnor \mul_19_13_g22610/U$1 ( \3893 , \3890 , \3892 );
mxor \mul_19_13_g22918/U$1 ( \3894 , \c[15] , \c[14] );
mxor \mul_19_13_g22874/U$1 ( \3895 , \b[0] , \c[15] );
mnand \mul_19_13_g22769/U$1 ( \3896 , \3894 , \3895 );
mor \mul_19_13_g22596/U$2 ( \3897 , \3896 , \2534 );
mxor \mul_19_13_g22889/U$1 ( \3898 , \b[1] , \c[15] );
mnand \mul_19_13_g22709/U$1 ( \3899 , \2534 , \3898 );
mnand \mul_19_13_g22596/U$1 ( \3900 , \3897 , \3899 );
mxor \g37115/U$1 ( \3901 , \3893 , \3900 );
mnot \mul_19_13_g22636/U$3 ( \3902 , \2505 );
mnot \mul_19_13_g22636/U$4 ( \3903 , \1743 );
mor \mul_19_13_g22636/U$2 ( \3904 , \3902 , \3903 );
mnot \mul_19_13_g22962/U$2 ( \3905 , \c[7] );
mnand \mul_19_13_g22962/U$1 ( \3906 , \3905 , \b[9] );
mnot \mul_19_13_g22714/U$3 ( \3907 , \3906 );
mnot \mul_19_13_g23078/U$2 ( \3908 , \b[9] );
mnand \mul_19_13_g23078/U$1 ( \3909 , \3908 , \c[7] );
mnot \mul_19_13_g22714/U$4 ( \3910 , \3909 );
mor \mul_19_13_g22714/U$2 ( \3911 , \3907 , \3910 );
mnand \mul_19_13_g22714/U$1 ( \3912 , \3911 , \1747 );
mnand \mul_19_13_g22636/U$1 ( \3913 , \3904 , \3912 );
mxnor \g37115/U$1_r1 ( \3914 , \3901 , \3913 );
mnot \mul_19_13_g37293/U$2 ( \3915 , \3914 );
mxor \mul_19_13_g37293/U$1 ( \3916 , \3889 , \3915 );
mxnor \g37113/U$1_r1 ( \3917 , \3885 , \3916 );
mxnor \mul_19_13_g23042/U$1 ( \3918 , \3859 , \3917 );
mxor \mul_19_13_g36760/U$1 ( \3919 , \3852 , \3918 );
mxnor \mul_19_13_g23036/U$1 ( \3920 , \3810 , \3919 );
mnot \mul_19_13_g22254/U$1 ( \3921 , \3920 );
mand \mul_19_13_g22231/U$2 ( \3922 , \3802 , \3921 );
mnot \mul_19_13_g22231/U$4 ( \3923 , \3802 );
mand \mul_19_13_g22231/U$3 ( \3924 , \3923 , \3920 );
mnor \mul_19_13_g22231/U$1 ( \3925 , \3922 , \3924 );
mnand \g4774/U$1 ( \3926 , \3925 , \2413 );
mnor \add_7_12_g9761/U$1 ( \3927 , \c[15] , \d[15] );
mnot \add_7_12_g9724/U$2 ( \3928 , \3927 );
mnand \add_7_12_g9752/U$1 ( \3929 , \c[15] , \d[15] );
mnand \add_7_12_g9724/U$1 ( \3930 , \3928 , \3929 );
mnand \add_7_12_g9741/U$1 ( \3931 , \c[1] , \d[1] );
mnand \add_7_12_g9770/U$1 ( \3932 , \c[0] , \d[0] );
mand \add_7_12_g9694/U$2 ( \3933 , \3931 , \3932 );
mnor \add_7_12_g9748/U$1 ( \3934 , \c[1] , \d[1] );
mnor \add_7_12_g9751/U$1 ( \3935 , \c[2] , \d[2] );
mnor \add_7_12_g9694/U$1 ( \3936 , \3933 , \3934 , \3935 );
mnot \add_7_12_g9775/U$2 ( \3937 , \3936 );
mnand \add_7_12_g9745/U$1 ( \3938 , \c[3] , \d[3] );
mnand \add_7_12_g9735/U$1 ( \3939 , \c[2] , \d[2] );
mnand \add_7_12_g9775/U$1 ( \3940 , \3937 , \3938 , \3939 );
mnor \add_7_12_g9746/U$1 ( \3941 , \c[5] , \d[5] );
mnor \add_7_12_g9755/U$1 ( \3942 , \c[4] , \d[4] );
mnor \add_7_12_g9727/U$1 ( \3943 , \3941 , \3942 );
mnor \add_7_12_g9739/U$1 ( \3944 , \c[7] , \d[7] );
mnor \add_7_12_g9737/U$1 ( \3945 , \c[6] , \d[6] );
mnor \add_7_12_g9732/U$1 ( \3946 , \3944 , \3945 );
mnor \add_7_12_g9754/U$1 ( \3947 , \c[3] , \d[3] );
mnot \add_7_12_g9753/U$1 ( \3948 , \3947 );
mnand \add_7_12_g9679/U$1 ( \3949 , \3940 , \3943 , \3946 , \3948 );
mnand \add_7_12_g9757/U$1 ( \3950 , \c[4] , \d[4] );
mnor \add_7_12_g9709/U$1 ( \3951 , \3941 , \3950 );
mnand \add_7_12_g9747/U$1 ( \3952 , \c[6] , \d[6] );
mnand \add_7_12_g9750/U$1 ( \3953 , \c[7] , \d[7] );
mnand \add_7_12_g9763/U$1 ( \3954 , \c[5] , \d[5] );
mnand \add_7_12_g9708/U$1 ( \3955 , \3952 , \3953 , \3954 );
mor \add_7_12_g9690/U$2 ( \3956 , \3951 , \3955 );
mnot \add_7_12_g9749/U$1 ( \3957 , \3953 );
mor \add_7_12_g9690/U$3 ( \3958 , \3946 , \3957 );
mnand \add_7_12_g9690/U$1 ( \3959 , \3956 , \3958 );
mnand \add_7_12_g9673/U$1 ( \3960 , \3949 , \3959 );
mnor \add_7_12_g9740/U$1 ( \3961 , \c[11] , \d[11] );
mnor \add_7_12_g9760/U$1 ( \3962 , \c[10] , \d[10] );
mnor \add_7_12_g9721/U$1 ( \3963 , \3961 , \3962 );
mnor \add_7_12_g9743/U$1 ( \3964 , \c[9] , \d[9] );
mnor \add_7_12_g9767/U$1 ( \3965 , \c[8] , \d[8] );
mnor \add_7_12_g9725/U$1 ( \3966 , \3964 , \3965 );
mnand \add_7_12_g9698/U$1 ( \3967 , \3963 , \3966 );
mnot \add_7_12_g9697/U$1 ( \3968 , \3967 );
mnor \add_7_12_g9769/U$1 ( \3969 , \c[14] , \d[14] );
mnot \add_7_12_g9700/U$2 ( \3970 , \3969 );
mnor \add_7_12_g9768/U$1 ( \3971 , \c[13] , \d[13] );
mnor \add_7_12_g9765/U$1 ( \3972 , \c[12] , \d[12] );
mnor \add_7_12_g9726/U$1 ( \3973 , \3971 , \3972 );
mnand \add_7_12_g9700/U$1 ( \3974 , \3970 , \3973 );
mnot \add_7_12_g9699/U$1 ( \3975 , \3974 );
mand \add_7_12_g9663/U$2 ( \3976 , \3960 , \3968 , \3975 );
mnand \add_7_12_g9738/U$1 ( \3977 , \c[8] , \d[8] );
mor \add_7_12_g9706/U$2 ( \3978 , \3964 , \3977 );
mnand \add_7_12_g9758/U$1 ( \3979 , \c[9] , \d[9] );
mnand \add_7_12_g9706/U$1 ( \3980 , \3978 , \3979 );
mand \add_7_12_g9692/U$2 ( \3981 , \3963 , \3980 );
mnand \add_7_12_g9762/U$1 ( \3982 , \c[10] , \d[10] );
mor \add_7_12_g9707/U$2 ( \3983 , \3961 , \3982 );
mnand \add_7_12_g9756/U$1 ( \3984 , \c[11] , \d[11] );
mnand \add_7_12_g9707/U$1 ( \3985 , \3983 , \3984 );
mnor \add_7_12_g9692/U$1 ( \3986 , \3981 , \3985 );
mor \add_7_12_g9682/U$2 ( \3987 , \3986 , \3974 );
mnand \add_7_12_g9742/U$1 ( \3988 , \c[12] , \d[12] );
mor \add_7_12_g9703/U$2 ( \3989 , \3971 , \3988 );
mnand \add_7_12_g9744/U$1 ( \3990 , \c[13] , \d[13] );
mnand \add_7_12_g9703/U$1 ( \3991 , \3989 , \3990 );
mnot \add_7_12_g9702/U$1 ( \3992 , \3991 );
mor \add_7_12_g9682/U$3 ( \3993 , \3969 , \3992 );
mnand \add_7_12_g9766/U$1 ( \3994 , \c[14] , \d[14] );
mnand \add_7_12_g9682/U$1 ( \3995 , \3987 , \3993 , \3994 );
mnor \add_7_12_g9663/U$1 ( \3996 , \3976 , \3995 );
mxor \add_7_12_g9646/U$1 ( \3997 , \3930 , \3996 );
mnot \add_7_12_g9719/U$2 ( \3998 , \3944 );
mnand \add_7_12_g9719/U$1 ( \3999 , \3998 , \3953 );
mor \add_7_12_g9688/U$2 ( \4000 , \3934 , \3932 );
mnand \add_7_12_g9688/U$1 ( \4001 , \4000 , \3931 );
mnor \add_7_12_g9716/U$1 ( \4002 , \3947 , \3935 );
mand \add_7_12_g9678/U$2 ( \4003 , \4001 , \4002 );
mor \add_7_12_g9704/U$2 ( \4004 , \3947 , \3939 );
mnand \add_7_12_g9704/U$1 ( \4005 , \4004 , \3938 );
mnor \add_7_12_g9678/U$1 ( \4006 , \4003 , \4005 );
mnot \add_7_12_g9677/U$1 ( \4007 , \4006 );
mnot \add_7_12_g9736/U$1 ( \4008 , \3945 );
mand \add_7_12_g9669/U$2 ( \4009 , \4007 , \3943 , \4008 );
mnot \add_7_12_g9687/U$3 ( \4010 , \4008 );
mnot \add_7_12_g9696/U$2 ( \4011 , \3951 );
mnand \add_7_12_g9696/U$1 ( \4012 , \4011 , \3954 );
mnot \add_7_12_g9687/U$4 ( \4013 , \4012 );
mor \add_7_12_g9687/U$2 ( \4014 , \4010 , \4013 );
mnand \add_7_12_g9687/U$1 ( \4015 , \4014 , \3952 );
mnor \add_7_12_g9669/U$1 ( \4016 , \4009 , \4015 );
mxor \add_7_12_g9653/U$1 ( \4017 , \3999 , \4016 );
mnand \add_7_12_g9720/U$1 ( \4018 , \4008 , \3952 );
mand \add_7_12_g9670/U$2 ( \4019 , \4007 , \3943 );
mnor \add_7_12_g9670/U$1 ( \4020 , \4019 , \4012 );
mxor \add_7_12_g9654/U$1 ( \4021 , \4018 , \4020 );
mnot \add_7_12_g9712/U$2 ( \4022 , \3954 );
mnor \add_7_12_g9712/U$1 ( \4023 , \4022 , \3941 );
mor \add_7_12_g9668/U$2 ( \4024 , \4006 , \3942 );
mnand \add_7_12_g9668/U$1 ( \4025 , \4024 , \3950 );
mxor \add_7_12_g9655/U$1 ( \4026 , \4023 , \4025 );
mand \add_7_12_g9657/U$2 ( \4027 , \3960 , \3966 );
mnor \add_7_12_g9657/U$1 ( \4028 , \4027 , \3980 );
mnot \add_7_12_g9764/U$1 ( \4029 , \3972 );
mand \add_7_12_g9659/U$2 ( \4030 , \3960 , \3968 , \4029 );
mor \add_7_12_g9676/U$2 ( \4031 , \3986 , \3972 );
mnand \add_7_12_g9676/U$1 ( \4032 , \4031 , \3988 );
mnor \add_7_12_g9659/U$1 ( \4033 , \4030 , \4032 );
mand \add_7_12_g9660/U$2 ( \4034 , \3960 , \3968 , \3973 );
mnot \add_7_12_g9675/U$2 ( \4035 , \3991 );
mnot \add_7_12_g9774/U$2 ( \4036 , \3986 );
mnand \add_7_12_g9774/U$1 ( \4037 , \4036 , \3973 );
mnand \add_7_12_g9675/U$1 ( \4038 , \4035 , \4037 );
mnor \add_7_12_g9660/U$1 ( \4039 , \4034 , \4038 );
mnot \add_7_12_g9672/U$1 ( \4040 , \3960 );
mor \add_7_12_g9662/U$2 ( \4041 , \4040 , \3965 );
mnand \add_7_12_g9662/U$1 ( \4042 , \4041 , \3977 );
mnor \add_7_12_g9728/U$1 ( \4043 , \3969 , \3927 );
mnand \add_7_12_g9701/U$1 ( \4044 , \4043 , \3973 );
mor \add_7_12_g9664/U$2 ( \4045 , \4040 , \3967 , \4044 );
mand \add_7_12_g9680/U$2 ( \4046 , \3991 , \4043 );
mnor \add_7_12_g9684/U$1 ( \4047 , \3986 , \4044 );
mor \add_7_12_g9705/U$2 ( \4048 , \3927 , \3994 );
mnand \add_7_12_g9705/U$1 ( \4049 , \4048 , \3929 );
mnor \add_7_12_g9680/U$1 ( \4050 , \4046 , \4047 , \4049 );
mnand \add_7_12_g9664/U$1 ( \4051 , \4045 , \4050 );
mnot \add_7_12_g9759/U$1 ( \4052 , \3962 );
mand \add_7_12_g9665/U$2 ( \4053 , \3960 , \3966 , \4052 );
mnot \add_7_12_g9689/U$3 ( \4054 , \4052 );
mnot \add_7_12_g9689/U$4 ( \4055 , \3980 );
mor \add_7_12_g9689/U$2 ( \4056 , \4054 , \4055 );
mnand \add_7_12_g9689/U$1 ( \4057 , \4056 , \3982 );
mnor \add_7_12_g9665/U$1 ( \4058 , \4053 , \4057 );
mor \add_7_12_g9666/U$2 ( \4059 , \4040 , \3967 );
mnand \add_7_12_g9666/U$1 ( \4060 , \4059 , \3986 );
mnot \add_7_12_g9718/U$2 ( \4061 , \3965 );
mnand \add_7_12_g9718/U$1 ( \4062 , \4061 , \3977 );
mand \add_7_12_g9667/U$2 ( \4063 , \4062 , \3960 );
mnot \add_7_12_g9667/U$4 ( \4064 , \4062 );
mand \add_7_12_g9667/U$3 ( \4065 , \4064 , \4040 );
mor \add_7_12_g9667/U$1 ( \4066 , \4063 , \4065 );
mnot \add_7_12_g9722/U$2 ( \4067 , \3942 );
mnand \add_7_12_g9722/U$1 ( \4068 , \4067 , \3950 );
mand \add_7_12_g9671/U$2 ( \4069 , \4068 , \4007 );
mnot \add_7_12_g9671/U$4 ( \4070 , \4068 );
mand \add_7_12_g9671/U$3 ( \4071 , \4070 , \4006 );
mor \add_7_12_g9671/U$1 ( \4072 , \4069 , \4071 );
mnand \add_7_12_g9731/U$1 ( \4073 , \3948 , \3938 );
mnot \add_7_12_g9683/U$2 ( \4074 , \3939 );
mnor \add_7_12_g9683/U$1 ( \4075 , \4074 , \3936 );
mxor \add_7_12_g9674/U$1 ( \4076 , \4073 , \4075 );
mnot \add_7_12_g9723/U$2 ( \4077 , \3939 );
mnor \add_7_12_g9723/U$1 ( \4078 , \4077 , \3935 );
mxor \add_7_12_g9681/U$1 ( \4079 , \4078 , \4001 );
mnot \add_7_12_g9729/U$2 ( \4080 , \3934 );
mnand \add_7_12_g9729/U$1 ( \4081 , \4080 , \3931 );
mxor \add_7_12_g9695/U$1 ( \4082 , \3932 , \4081 );
mnand \add_7_12_g9711/U$1 ( \4083 , \4029 , \3988 );
mnot \add_7_12_g9714/U$2 ( \4084 , \3961 );
mnand \add_7_12_g9714/U$1 ( \4085 , \4084 , \3984 );
mnand \add_7_12_g9715/U$1 ( \4086 , \4052 , \3982 );
mnot \add_7_12_g9717/U$2 ( \4087 , \3979 );
mnor \add_7_12_g9717/U$1 ( \4088 , \4087 , \3964 );
mnot \add_7_12_g9730/U$2 ( \4089 , \3969 );
mnand \add_7_12_g9730/U$1 ( \4090 , \4089 , \3994 );
mnot \add_7_12_g9733/U$2 ( \4091 , \3971 );
mnand \add_7_12_g9733/U$1 ( \4092 , \4091 , \3990 );
mxor \add_7_12_g2/U$1 ( \4093 , \4086 , \4028 );
mxor \add_7_12_g9772/U$1 ( \4094 , \4092 , \4033 );
mxor \add_7_12_g9773/U$1 ( \4095 , \4088 , \4042 );
mxnor \add_7_12_g9776/U$1 ( \4096 , \4060 , \4083 );
mxor \add_7_12_g9777/U$1 ( \4097 , \4058 , \4085 );
mxor \add_7_12_g9778/U$1 ( \4098 , \d[0] , \c[0] );
mnand \g36996/U$1 ( \4099 , \3926 , \3788 , \3517 , \927 );
mbuf \mul_7_15_fopt36211/U$1 ( \4100 , \4099 );
mnot \mul_7_15_fopt36210/U$1 ( \4101 , \4100 );
mnot \mul_7_15_fopt36207/U$1 ( \4102 , \4101 );
mand \mul_7_15_g35783/U$1 ( \4103 , \4102 , \4096 );
mnot \mul_7_15_g35679/U$3 ( \4104 , \3997 );
mbuf \fopt36879/U$1 ( \4105 , \2477 );
mbuf \fopt36878/U$1 ( \4106 , \4105 );
mnot \fopt36874/U$1 ( \4107 , \4106 );
mnot \mul_7_15_g35679/U$4 ( \4108 , \4107 );
mor \mul_7_15_g35679/U$2 ( \4109 , \4104 , \4108 );
mbuf \fopt36862/U$1 ( \4110 , \4105 );
mnot \mul_7_15_g36081/U$1 ( \4111 , \3997 );
mnand \mul_7_15_g35819/U$1 ( \4112 , \4110 , \4111 );
mnand \mul_7_15_g35679/U$1 ( \4113 , \4109 , \4112 );
mnot \mul_7_15_g35135/U$3 ( \4114 , \4113 );
mnand \g37035/U$1 ( \4115 , \3193 , \3656 );
mnot \mul_7_15_g36019/U$1 ( \4116 , \4115 );
mnot \mul_7_15_g35563/U$3 ( \4117 , \4116 );
mnot \mul_7_15_g35563/U$4 ( \4118 , \4105 );
mor \mul_7_15_g35563/U$2 ( \4119 , \4117 , \4118 );
mnot \g37102/U$3 ( \4120 , \3656 );
mnot \g37102/U$4 ( \4121 , \3193 );
mor \g37102/U$2 ( \4122 , \4120 , \4121 );
mnot \fopt36863/U$1 ( \4123 , \4105 );
mnand \g37102/U$1 ( \4124 , \4122 , \4123 );
mnand \mul_7_15_g35563/U$1 ( \4125 , \4119 , \4124 );
mxnor \g36553/U$1 ( \4126 , \2876 , \4115 );
mnand \mul_7_15_g35459/U$1 ( \4127 , \4125 , \4126 );
mnot \mul_7_15_g35458/U$1 ( \4128 , \4127 );
mbuf \mul_7_15_g35456_dup/U$1 ( \4129 , \4128 );
mnot \mul_7_15_g35135/U$4 ( \4130 , \4129 );
mor \mul_7_15_g35135/U$2 ( \4131 , \4114 , \4130 );
mnot \mul_7_15_g35561/U$1 ( \4132 , \4126 );
mbuf \mul_7_15_g35557/U$1 ( \4133 , \4132 );
mnot \fopt36861/U$1 ( \4134 , \4110 );
mnot \mul_7_15_g36080/U$1 ( \4135 , \4051 );
mand \g37077/U$2 ( \4136 , \4134 , \4135 );
mnot \g37077/U$4 ( \4137 , \4134 );
mand \g37077/U$3 ( \4138 , \4137 , \4051 );
mnor \g37077/U$1 ( \4139 , \4136 , \4138 );
mnand \mul_7_15_g35364/U$1 ( \4140 , \4133 , \4139 );
mnand \mul_7_15_g35135/U$1 ( \4141 , \4131 , \4140 );
mxor \mul_7_15_g34814/U$1 ( \4142 , \4103 , \4141 );
mnot \fopt36787/U$1 ( \4143 , \3637 );
mnot \mul_7_15_g35570/U$3 ( \4144 , \4143 );
mnot \mul_7_15_g35570/U$4 ( \4145 , \3573 );
mor \mul_7_15_g35570/U$2 ( \4146 , \4144 , \4145 );
mnot \mul_7_15_fopt36217/U$1 ( \4147 , \3573 );
mnand \mul_7_15_g35759/U$1 ( \4148 , \4147 , \3637 );
mnand \mul_7_15_g35570/U$1 ( \4149 , \4146 , \4148 );
mbuf \mul_7_15_g35569/U$1 ( \4150 , \4149 );
mnot \mul_7_15_g35568/U$1 ( \4151 , \4150 );
mnot \mul_7_15_g35028/U$3 ( \4152 , \4151 );
mnot \mul_7_15_g36047/U$1 ( \4153 , \2876 );
mnot \mul_7_15_g36028/U$1 ( \4154 , \4153 );
mand \mul_7_15_g35571/U$2 ( \4155 , \4154 , \4147 );
mand \mul_7_15_g35571/U$3 ( \4156 , \4153 , \3573 );
mnor \mul_7_15_g35571/U$1 ( \4157 , \4155 , \4156 );
mnor \mul_7_15_g35415/U$1 ( \4158 , \4157 , \4149 );
mbuf \fopt36883/U$1 ( \4159 , \4158 );
mnot \fopt36884/U$1 ( \4160 , \4159 );
mnot \mul_7_15_g35028/U$4 ( \4161 , \4160 );
mor \mul_7_15_g35028/U$2 ( \4162 , \4152 , \4161 );
mbuf \mul_7_15_g36046/U$1 ( \4163 , \4153 );
mnot \mul_7_15_g36031/U$1 ( \4164 , \4163 );
mnand \mul_7_15_g35028/U$1 ( \4165 , \4162 , \4164 );
mxor \mul_7_15_g34814/U$1_r1 ( \4166 , \4142 , \4165 );
mnot \mul_7_15_g35614/U$3 ( \4167 , \4051 );
mnot \mul_7_15_g35614/U$4 ( \4168 , \4163 );
mor \mul_7_15_g35614/U$2 ( \4169 , \4167 , \4168 );
mnot \mul_7_15_g36033/U$1 ( \4170 , \4163 );
mnand \mul_7_15_g35791/U$1 ( \4171 , \4135 , \4170 );
mnand \mul_7_15_g35614/U$1 ( \4172 , \4169 , \4171 );
mnot \mul_7_15_g35246/U$3 ( \4173 , \4172 );
mnot \mul_7_15_g35246/U$4 ( \4174 , \4159 );
mor \mul_7_15_g35246/U$2 ( \4175 , \4173 , \4174 );
mnand \mul_7_15_g35487/U$1 ( \4176 , \4150 , \4164 );
mnand \mul_7_15_g35246/U$1 ( \4177 , \4175 , \4176 );
mxor \mul_7_15_g35511/U$1 ( \4178 , \4094 , \4100 );
mnot \mul_7_15_g35054/U$3 ( \4179 , \4178 );
mnot \fopt36966/U$1 ( \4180 , \2790 );
mnot \fopt36965/U$1 ( \4181 , \4180 );
mnot \fopt36963/U$1 ( \4182 , \4181 );
mnand \mul_7_15_g35763/U$1 ( \4183 , \4099 , \4182 );
mnot \mul_7_15_g35403/U$3 ( \4184 , \4183 );
mand \g36995/U$1 ( \4185 , \3926 , \3788 , \3517 , \927 );
mnand \mul_7_15_g35761/U$1 ( \4186 , \4181 , \4185 );
mnot \mul_7_15_g35403/U$4 ( \4187 , \4186 );
mor \mul_7_15_g35403/U$2 ( \4188 , \4184 , \4187 );
mand \mul_7_15_g35541/U$2 ( \4189 , \2477 , \2790 );
mnot \mul_7_15_g35541/U$4 ( \4190 , \2477 );
mand \mul_7_15_g35541/U$3 ( \4191 , \4190 , \4180 );
mor \mul_7_15_g35541/U$1 ( \4192 , \4189 , \4191 );
mnand \mul_7_15_g35403/U$1 ( \4193 , \4188 , \4192 );
mnot \fopt36855/U$1 ( \4194 , \4193 );
mbuf \fopt36854/U$1 ( \4195 , \4194 );
mnot \mul_7_15_g35054/U$4 ( \4196 , \4195 );
mor \mul_7_15_g35054/U$2 ( \4197 , \4179 , \4196 );
mxor \add_7_12_g37294/U$1 ( \4198 , \4039 , \4090 );
mxor \mul_7_15_g35516/U$1 ( \4199 , \4198 , \4102 );
mnot \mul_7_15_g35540/U$1 ( \4200 , \4192 );
mnand \mul_7_15_g35255/U$1 ( \4201 , \4199 , \4200 );
mnand \mul_7_15_g35054/U$1 ( \4202 , \4197 , \4201 );
mxor \mul_7_15_g34670/U$1 ( \4203 , \4177 , \4202 );
mand \mul_7_15_g35782/U$1 ( \4204 , \4102 , \4097 );
mnot \mul_7_15_g35648/U$3 ( \4205 , \4198 );
mnot \fopt36871/U$1 ( \4206 , \4106 );
mnot \mul_7_15_g35648/U$4 ( \4207 , \4206 );
mor \mul_7_15_g35648/U$2 ( \4208 , \4205 , \4207 );
mnot \mul_7_15_g35944/U$1 ( \4209 , \4198 );
mnand \mul_7_15_g35852/U$1 ( \4210 , \4110 , \4209 );
mnand \mul_7_15_g35648/U$1 ( \4211 , \4208 , \4210 );
mnot \mul_7_15_g35167/U$3 ( \4212 , \4211 );
mnot \mul_7_15_g35167/U$4 ( \4213 , \4129 );
mor \mul_7_15_g35167/U$2 ( \4214 , \4212 , \4213 );
mnand \mul_7_15_g35387/U$1 ( \4215 , \4133 , \4113 );
mnand \mul_7_15_g35167/U$1 ( \4216 , \4214 , \4215 );
mxor \mul_7_15_g34752/U$4 ( \4217 , \4204 , \4216 );
mand \mul_7_15_g35600/U$2 ( \4218 , \4096 , \4100 );
mnot \mul_7_15_g35600/U$4 ( \4219 , \4096 );
mand \mul_7_15_g35600/U$3 ( \4220 , \4219 , \4101 );
mnor \mul_7_15_g35600/U$1 ( \4221 , \4218 , \4220 );
mnot \mul_7_15_g35060/U$3 ( \4222 , \4221 );
mnot \mul_7_15_g35060/U$4 ( \4223 , \4195 );
mor \mul_7_15_g35060/U$2 ( \4224 , \4222 , \4223 );
mnand \mul_7_15_g35249/U$1 ( \4225 , \4178 , \4200 );
mnand \mul_7_15_g35060/U$1 ( \4226 , \4224 , \4225 );
mand \mul_7_15_g34752/U$3 ( \4227 , \4217 , \4226 );
mand \mul_7_15_g34752/U$5 ( \4228 , \4204 , \4216 );
mor \mul_7_15_g34752/U$2 ( \4229 , \4227 , \4228 );
mxor \mul_7_15_g34670/U$1_r1 ( \4230 , \4203 , \4229 );
mxor \mul_7_15_g34517/U$1 ( \4231 , \4166 , \4230 );
mnot \mul_7_15_g34679/U$3 ( \4232 , \4177 );
mxor \mul_7_15_g34752/U$1 ( \4233 , \4204 , \4216 );
mxor \mul_7_15_g34752/U$1_r1 ( \4234 , \4233 , \4226 );
mnot \mul_7_15_g34750/U$1 ( \4235 , \4234 );
mnot \mul_7_15_g34679/U$4 ( \4236 , \4235 );
mor \mul_7_15_g34679/U$2 ( \4237 , \4232 , \4236 );
mnot \mul_7_15_g35623/U$3 ( \4238 , \3997 );
mnot \mul_7_15_g35623/U$4 ( \4239 , \4163 );
mor \mul_7_15_g35623/U$2 ( \4240 , \4238 , \4239 );
mnand \mul_7_15_g35796/U$1 ( \4241 , \4170 , \4111 );
mnand \mul_7_15_g35623/U$1 ( \4242 , \4240 , \4241 );
mnot \mul_7_15_g35171/U$3 ( \4243 , \4242 );
mnot \mul_7_15_g35171/U$4 ( \4244 , \4159 );
mor \mul_7_15_g35171/U$2 ( \4245 , \4243 , \4244 );
mnand \mul_7_15_g35416/U$1 ( \4246 , \4150 , \4172 );
mnand \mul_7_15_g35171/U$1 ( \4247 , \4245 , \4246 );
mnot \mul_7_15_g34905/U$3 ( \4248 , \4247 );
mnot \mul_7_15_g35610/U$3 ( \4249 , \4097 );
mnot \mul_7_15_fopt36196/U$1 ( \4250 , \4100 );
mnot \mul_7_15_g35610/U$4 ( \4251 , \4250 );
mor \mul_7_15_g35610/U$2 ( \4252 , \4249 , \4251 );
mnot \mul_7_15_fopt36199/U$1 ( \4253 , \4101 );
mnot \mul_7_15_g36023/U$1 ( \4254 , \4097 );
mnand \mul_7_15_g35830/U$1 ( \4255 , \4253 , \4254 );
mnand \mul_7_15_g35610/U$1 ( \4256 , \4252 , \4255 );
mnot \mul_7_15_g35066/U$3 ( \4257 , \4256 );
mnot \mul_7_15_g35066/U$4 ( \4258 , \4195 );
mor \mul_7_15_g35066/U$2 ( \4259 , \4257 , \4258 );
mnand \mul_7_15_g35256/U$1 ( \4260 , \4221 , \4200 );
mnand \mul_7_15_g35066/U$1 ( \4261 , \4259 , \4260 );
mnot \mul_7_15_g34905/U$4 ( \4262 , \4261 );
mor \mul_7_15_g34905/U$2 ( \4263 , \4248 , \4262 );
mor \mul_7_15_g34943/U$2 ( \4264 , \4261 , \4247 );
mxnor \mul_7_15_g36433/U$1 ( \4265 , \3136 , \3326 );
mnot \mul_7_15_g35582/U$1 ( \4266 , \4265 );
mnot \mul_7_15_g35581/U$1 ( \4267 , \4266 );
mbuf \mul_7_15_g35580/U$1 ( \4268 , \4267 );
mnot \mul_7_15_g35030/U$3 ( \4269 , \4268 );
mnot \mul_7_15_g35917/U$1 ( \4270 , \3136 );
mnand \mul_7_15_g35769/U$1 ( \4271 , \4270 , \3637 );
mnot \mul_7_15_g35315/U$3 ( \4272 , \4271 );
mnot \mul_7_15_g36435/U$2 ( \4273 , \3637 );
mnot \mul_7_15_g35916/U$1 ( \4274 , \4270 );
mnand \mul_7_15_g36435/U$1 ( \4275 , \4273 , \4274 );
mnot \mul_7_15_g35315/U$4 ( \4276 , \4275 );
mor \mul_7_15_g35315/U$2 ( \4277 , \4272 , \4276 );
mnand \mul_7_15_g35315/U$1 ( \4278 , \4277 , \4265 );
mnot \fopt36701/U$1 ( \4279 , \4278 );
mnot \fopt36699/U$1 ( \4280 , \4279 );
mnot \mul_7_15_g35030/U$4 ( \4281 , \4280 );
mor \mul_7_15_g35030/U$2 ( \4282 , \4269 , \4281 );
mbuf \fopt36804/U$1 ( \4283 , \3637 );
mnot \fopt36803/U$1 ( \4284 , \4283 );
mnot \fopt36801/U$1 ( \4285 , \4284 );
mnand \mul_7_15_g35030/U$1 ( \4286 , \4282 , \4285 );
mnand \mul_7_15_g34943/U$1 ( \4287 , \4264 , \4286 );
mnand \mul_7_15_g34905/U$1 ( \4288 , \4263 , \4287 );
mnand \mul_7_15_g34679/U$1 ( \4289 , \4237 , \4288 );
mnot \mul_7_15_g36418/U$2 ( \4290 , \4177 );
mnand \mul_7_15_g36418/U$1 ( \4291 , \4290 , \4234 );
mnand \mul_7_15_g34655/U$1 ( \4292 , \4289 , \4291 );
mxnor \mul_7_15_g34517/U$1_r1 ( \4293 , \4231 , \4292 );
mand \mul_7_15_g35775/U$1 ( \4294 , \4102 , \4093 );
mnot \mul_7_15_g35639/U$3 ( \4295 , \4094 );
mnot \mul_7_15_g35639/U$4 ( \4296 , \4206 );
mor \mul_7_15_g35639/U$2 ( \4297 , \4295 , \4296 );
mnot \mul_7_15_g36022/U$1 ( \4298 , \4094 );
mnand \mul_7_15_g35836/U$1 ( \4299 , \4106 , \4298 );
mnand \mul_7_15_g35639/U$1 ( \4300 , \4297 , \4299 );
mnot \mul_7_15_g35180/U$3 ( \4301 , \4300 );
mbuf \mul_7_15_g36999/U$1 ( \4302 , \4128 );
mnot \mul_7_15_g35180/U$4 ( \4303 , \4302 );
mor \mul_7_15_g35180/U$2 ( \4304 , \4301 , \4303 );
mnand \mul_7_15_g35428/U$1 ( \4305 , \4133 , \4211 );
mnand \mul_7_15_g35180/U$1 ( \4306 , \4304 , \4305 );
mxor \mul_7_15_g34773/U$4 ( \4307 , \4294 , \4306 );
mnot \mul_7_15_g35649/U$3 ( \4308 , \4198 );
mnot \mul_7_15_g35649/U$4 ( \4309 , \4163 );
mor \mul_7_15_g35649/U$2 ( \4310 , \4308 , \4309 );
mnot \mul_7_15_g36036/U$1 ( \4311 , \4163 );
mnand \mul_7_15_g35858/U$1 ( \4312 , \4311 , \4209 );
mnand \mul_7_15_g35649/U$1 ( \4313 , \4310 , \4312 );
mnot \mul_7_15_g35203/U$3 ( \4314 , \4313 );
mnot \mul_7_15_g35203/U$4 ( \4315 , \4159 );
mor \mul_7_15_g35203/U$2 ( \4316 , \4314 , \4315 );
mbuf \mul_7_15_g35564/U$1 ( \4317 , \4150 );
mnand \mul_7_15_g35337/U$1 ( \4318 , \4317 , \4242 );
mnand \mul_7_15_g35203/U$1 ( \4319 , \4316 , \4318 );
mand \mul_7_15_g34773/U$3 ( \4320 , \4307 , \4319 );
mand \mul_7_15_g34773/U$5 ( \4321 , \4294 , \4306 );
mor \mul_7_15_g34773/U$2 ( \4322 , \4320 , \4321 );
mnot \mul_7_15_g34574/U$2 ( \4323 , \4322 );
mxor \mul_7_15_g34658/U$1 ( \4324 , \4177 , \4288 );
mxnor \mul_7_15_g34658/U$1_r1 ( \4325 , \4324 , \4234 );
mnot \mul_7_15_g34634/U$1 ( \4326 , \4325 );
mnand \mul_7_15_g34574/U$1 ( \4327 , \4323 , \4326 );
mxor \mul_7_15_g34773/U$1 ( \4328 , \4294 , \4306 );
mxor \mul_7_15_g34773/U$1_r1 ( \4329 , \4328 , \4319 );
mand \mul_7_15_g35780/U$1 ( \4330 , \4102 , \4095 );
mnot \mul_7_15_g35615/U$3 ( \4331 , \4051 );
mnot \fopt36791/U$1 ( \4332 , \3637 );
mnot \mul_7_15_g35615/U$4 ( \4333 , \4332 );
mor \mul_7_15_g35615/U$2 ( \4334 , \4331 , \4333 );
mnand \mul_7_15_g35790/U$1 ( \4335 , \4283 , \4135 );
mnand \mul_7_15_g35615/U$1 ( \4336 , \4334 , \4335 );
mnot \mul_7_15_g35240/U$3 ( \4337 , \4336 );
mnot \fopt36697/U$1 ( \4338 , \4280 );
mnot \mul_7_15_g35240/U$4 ( \4339 , \4338 );
mor \mul_7_15_g35240/U$2 ( \4340 , \4337 , \4339 );
mnot \mul_7_15_g35579/U$1 ( \4341 , \4268 );
mnand \mul_7_15_g35488/U$1 ( \4342 , \4341 , \4285 );
mnand \mul_7_15_g35240/U$1 ( \4343 , \4340 , \4342 );
mxor \mul_7_15_g34774/U$4 ( \4344 , \4330 , \4343 );
mnot \mul_7_15_g35608/U$3 ( \4345 , \4093 );
mnot \mul_7_15_fopt36190/U$1 ( \4346 , \4100 );
mnot \mul_7_15_g35608/U$4 ( \4347 , \4346 );
mor \mul_7_15_g35608/U$2 ( \4348 , \4345 , \4347 );
mnot \mul_7_15_g36025/U$1 ( \4349 , \4093 );
mnand \mul_7_15_g35854/U$1 ( \4350 , \4100 , \4349 );
mnand \mul_7_15_g35608/U$1 ( \4351 , \4348 , \4350 );
mnot \mul_7_15_g35056/U$3 ( \4352 , \4351 );
mnot \mul_7_15_g35056/U$4 ( \4353 , \4195 );
mor \mul_7_15_g35056/U$2 ( \4354 , \4352 , \4353 );
mnand \mul_7_15_g35263/U$1 ( \4355 , \4256 , \4200 );
mnand \mul_7_15_g35056/U$1 ( \4356 , \4354 , \4355 );
mand \mul_7_15_g34774/U$3 ( \4357 , \4344 , \4356 );
mand \mul_7_15_g34774/U$5 ( \4358 , \4330 , \4343 );
mor \mul_7_15_g34774/U$2 ( \4359 , \4357 , \4358 );
mxor \mul_7_15_g34592/U$4 ( \4360 , \4329 , \4359 );
mxor \g37295/U$1 ( \4361 , \4286 , \4247 );
mxor \g37295/U$1_r1 ( \4362 , \4361 , \4261 );
mand \mul_7_15_g34592/U$3 ( \4363 , \4360 , \4362 );
mand \mul_7_15_g34592/U$5 ( \4364 , \4329 , \4359 );
mor \mul_7_15_g34592/U$2 ( \4365 , \4363 , \4364 );
mand \mul_7_15_g34491/U$2 ( \4366 , \4327 , \4365 );
mnot \mul_7_15_g36386/U$2 ( \4367 , \4322 );
mnor \mul_7_15_g36386/U$1 ( \4368 , \4367 , \4326 );
mnor \mul_7_15_g34491/U$1 ( \4369 , \4366 , \4368 );
mnand \mul_7_15_g34440/U$1 ( \4370 , \4293 , \4369 );
mnot \mul_7_15_g36367/U$2 ( \4371 , \4370 );
mnot \mul_7_15_g35945/U$1 ( \4372 , \4096 );
mnot \mul_7_15_g35668/U$3 ( \4373 , \4372 );
mnot \mul_7_15_g35668/U$4 ( \4374 , \4106 );
mor \mul_7_15_g35668/U$2 ( \4375 , \4373 , \4374 );
mnand \mul_7_15_g35889/U$1 ( \4376 , \4206 , \4096 );
mnand \mul_7_15_g35668/U$1 ( \4377 , \4375 , \4376 );
mnot \mul_7_15_g35214/U$3 ( \4378 , \4377 );
mnot \mul_7_15_g35214/U$4 ( \4379 , \4302 );
mor \mul_7_15_g35214/U$2 ( \4380 , \4378 , \4379 );
mnand \mul_7_15_g35346/U$1 ( \4381 , \4133 , \4300 );
mnand \mul_7_15_g35214/U$1 ( \4382 , \4380 , \4381 );
mnot \mul_7_15_g36415/U$2 ( \4383 , \4382 );
mnand \mul_7_15_g36415/U$1 ( \4384 , \4383 , \4319 );
mnot \mul_7_15_g34724/U$3 ( \4385 , \4384 );
mand \mul_7_15_g35772/U$1 ( \4386 , \4100 , \4066 );
mnot \mul_7_15_g35603/U$3 ( \4387 , \4095 );
mnot \mul_7_15_fopt36192/U$1 ( \4388 , \4100 );
mnot \mul_7_15_g35603/U$4 ( \4389 , \4388 );
mor \mul_7_15_g35603/U$2 ( \4390 , \4387 , \4389 );
mnot \mul_7_15_g36020/U$1 ( \4391 , \4095 );
mnand \mul_7_15_g35870/U$1 ( \4392 , \4100 , \4391 );
mnand \mul_7_15_g35603/U$1 ( \4393 , \4390 , \4392 );
mnot \mul_7_15_g35061/U$3 ( \4394 , \4393 );
mnot \fopt36849/U$1 ( \4395 , \4193 );
mnot \mul_7_15_g35061/U$4 ( \4396 , \4395 );
mor \mul_7_15_g35061/U$2 ( \4397 , \4394 , \4396 );
mnand \mul_7_15_g35254/U$1 ( \4398 , \4200 , \4351 );
mnand \mul_7_15_g35061/U$1 ( \4399 , \4397 , \4398 );
mxor \mul_7_15_g34831/U$4 ( \4400 , \4386 , \4399 );
mnot \mul_7_15_g35112/U$3 ( \4401 , \4159 );
mnot \mul_7_15_g35659/U$3 ( \4402 , \4094 );
mnot \mul_7_15_g35659/U$4 ( \4403 , \4163 );
mor \mul_7_15_g35659/U$2 ( \4404 , \4402 , \4403 );
mnand \mul_7_15_g35874/U$1 ( \4405 , \4170 , \4298 );
mnand \mul_7_15_g35659/U$1 ( \4406 , \4404 , \4405 );
mnot \mul_7_15_g35112/U$4 ( \4407 , \4406 );
mor \mul_7_15_g35112/U$2 ( \4408 , \4401 , \4407 );
mnand \mul_7_15_g35388/U$1 ( \4409 , \4150 , \4313 );
mnand \mul_7_15_g35112/U$1 ( \4410 , \4408 , \4409 );
mand \mul_7_15_g34831/U$3 ( \4411 , \4400 , \4410 );
mand \mul_7_15_g34831/U$5 ( \4412 , \4386 , \4399 );
mor \mul_7_15_g34831/U$2 ( \4413 , \4411 , \4412 );
mnot \mul_7_15_g34724/U$4 ( \4414 , \4413 );
mor \mul_7_15_g34724/U$2 ( \4415 , \4385 , \4414 );
mnot \mul_7_15_g36414/U$2 ( \4416 , \4319 );
mnand \mul_7_15_g36414/U$1 ( \4417 , \4416 , \4382 );
mnand \mul_7_15_g34724/U$1 ( \4418 , \4415 , \4417 );
mxor \mul_7_15_g34592/U$1 ( \4419 , \4329 , \4359 );
mxor \mul_7_15_g34592/U$1_r1 ( \4420 , \4419 , \4362 );
mxor \mul_7_15_g34452/U$1 ( \4421 , \4418 , \4420 );
mxor \mul_7_15_g34774/U$1 ( \4422 , \4330 , \4343 );
mxor \mul_7_15_g34774/U$1_r1 ( \4423 , \4422 , \4356 );
mnot \mul_7_15_g35626/U$3 ( \4424 , \3997 );
mnot \mul_7_15_g35626/U$4 ( \4425 , \4332 );
mor \mul_7_15_g35626/U$2 ( \4426 , \4424 , \4425 );
mnand \mul_7_15_g35802/U$1 ( \4427 , \4283 , \4111 );
mnand \mul_7_15_g35626/U$1 ( \4428 , \4426 , \4427 );
mnot \mul_7_15_g35147/U$3 ( \4429 , \4428 );
mbuf \fopt36700/U$1 ( \4430 , \4279 );
mnot \mul_7_15_g35147/U$4 ( \4431 , \4430 );
mor \mul_7_15_g35147/U$2 ( \4432 , \4429 , \4431 );
mnand \mul_7_15_g35344/U$1 ( \4433 , \4341 , \4336 );
mnand \mul_7_15_g35147/U$1 ( \4434 , \4432 , \4433 );
mnot \mul_7_15_fopt36243/U$1 ( \4435 , \3326 );
mnot \mul_7_15_fopt36242/U$1 ( \4436 , \4435 );
mnot \mul_7_15_g36015/U$1 ( \4437 , \3387 );
mand \mul_7_15_g35584/U$2 ( \4438 , \4436 , \4437 );
mand \mul_7_15_g35584/U$3 ( \4439 , \3387 , \4435 );
mnor \mul_7_15_g35584/U$1 ( \4440 , \4438 , \4439 );
mnot \mul_7_15_g35549/U$3 ( \4441 , \3387 );
mnot \mul_7_15_g36136/U$1 ( \4442 , \3448 );
mnot \mul_7_15_g35549/U$4 ( \4443 , \4442 );
mor \mul_7_15_g35549/U$2 ( \4444 , \4441 , \4443 );
mnot \mul_7_15_g36016/U$1 ( \4445 , \3387 );
mnand \mul_7_15_g35768/U$1 ( \4446 , \4445 , \3448 );
mnand \mul_7_15_g35549/U$1 ( \4447 , \4444 , \4446 );
mnor \mul_7_15_g35324/U$1 ( \4448 , \4440 , \4447 );
mbuf \mul_7_15_g35323/U$1 ( \4449 , \4448 );
mnot \mul_7_15_g35319/U$1 ( \4450 , \4449 );
mnot \mul_7_15_g35027/U$3 ( \4451 , \4450 );
mbuf \mul_7_15_g35548/U$1 ( \4452 , \4447 );
mbuf \mul_7_15_g35546/U$1 ( \4453 , \4452 );
mnot \mul_7_15_g35542/U$1 ( \4454 , \4453 );
mnot \mul_7_15_g35027/U$4 ( \4455 , \4454 );
mor \mul_7_15_g35027/U$2 ( \4456 , \4451 , \4455 );
mbuf \mul_7_15_fopt36230/U$1 ( \4457 , \4435 );
mnot \mul_7_15_fopt36218/U$1 ( \4458 , \4457 );
mnand \mul_7_15_g35027/U$1 ( \4459 , \4456 , \4458 );
mxor \mul_7_15_g34808/U$4 ( \4460 , \4434 , \4459 );
mand \mul_7_15_g35675/U$2 ( \4461 , \4097 , \4107 );
mnot \mul_7_15_g35675/U$4 ( \4462 , \4097 );
mand \mul_7_15_g35675/U$3 ( \4463 , \4462 , \4106 );
mnor \mul_7_15_g35675/U$1 ( \4464 , \4461 , \4463 );
mnot \mul_7_15_g35674/U$1 ( \4465 , \4464 );
mnot \mul_7_15_g35146/U$3 ( \4466 , \4465 );
mnot \mul_7_15_g35146/U$4 ( \4467 , \4129 );
mor \mul_7_15_g35146/U$2 ( \4468 , \4466 , \4467 );
mnand \mul_7_15_g35421/U$1 ( \4469 , \4133 , \4377 );
mnand \mul_7_15_g35146/U$1 ( \4470 , \4468 , \4469 );
mand \mul_7_15_g34808/U$3 ( \4471 , \4460 , \4470 );
mand \mul_7_15_g34808/U$5 ( \4472 , \4434 , \4459 );
mor \mul_7_15_g34808/U$2 ( \4473 , \4471 , \4472 );
mxor \mul_7_15_g34569/U$4 ( \4474 , \4423 , \4473 );
mnot \mul_7_15_g34946/U$3 ( \4475 , \4382 );
mnot \mul_7_15_g34946/U$4 ( \4476 , \4319 );
mand \mul_7_15_g34946/U$2 ( \4477 , \4475 , \4476 );
mand \mul_7_15_g34946/U$5 ( \4478 , \4382 , \4319 );
mnor \mul_7_15_g34946/U$1 ( \4479 , \4477 , \4478 );
mnot \mul_7_15_g34727/U$3 ( \4480 , \4479 );
mnot \mul_7_15_g34727/U$4 ( \4481 , \4413 );
mor \mul_7_15_g34727/U$2 ( \4482 , \4480 , \4481 );
mor \mul_7_15_g34727/U$5 ( \4483 , \4413 , \4479 );
mnand \mul_7_15_g34727/U$1 ( \4484 , \4482 , \4483 );
mand \mul_7_15_g34569/U$3 ( \4485 , \4474 , \4484 );
mand \mul_7_15_g34569/U$5 ( \4486 , \4423 , \4473 );
mor \mul_7_15_g34569/U$2 ( \4487 , \4485 , \4486 );
mxor \mul_7_15_g34452/U$1_r1 ( \4488 , \4421 , \4487 );
mnot \fopt36950/U$1 ( \4489 , \4488 );
mxor \mul_7_15_g34831/U$1 ( \4490 , \4386 , \4399 );
mxor \mul_7_15_g34831/U$1_r1 ( \4491 , \4490 , \4410 );
mnot \mul_7_15_g35697/U$3 ( \4492 , \4198 );
mnot \fopt36794/U$1 ( \4493 , \4283 );
mnot \mul_7_15_g35697/U$4 ( \4494 , \4493 );
mor \mul_7_15_g35697/U$2 ( \4495 , \4492 , \4494 );
mnand \mul_7_15_g35806/U$1 ( \4496 , \4285 , \4209 );
mnand \mul_7_15_g35697/U$1 ( \4497 , \4495 , \4496 );
mnot \mul_7_15_g35210/U$3 ( \4498 , \4497 );
mnot \mul_7_15_g35210/U$4 ( \4499 , \4338 );
mor \mul_7_15_g35210/U$2 ( \4500 , \4498 , \4499 );
mnand \mul_7_15_g35352/U$1 ( \4501 , \4341 , \4428 );
mnand \mul_7_15_g35210/U$1 ( \4502 , \4500 , \4501 );
mor \mul_7_15_g34719/U$2 ( \4503 , \4491 , \4502 );
mand \mul_7_15_g35633/U$2 ( \4504 , \4093 , \4134 );
mnot \mul_7_15_g35633/U$4 ( \4505 , \4093 );
mand \mul_7_15_g35633/U$3 ( \4506 , \4505 , \4106 );
mnor \mul_7_15_g35633/U$1 ( \4507 , \4504 , \4506 );
mnot \mul_7_15_g35173/U$3 ( \4508 , \4507 );
mnot \mul_7_15_g35173/U$4 ( \4509 , \4127 );
mand \mul_7_15_g35173/U$2 ( \4510 , \4508 , \4509 );
mnot \mul_7_15_g35560/U$1 ( \4511 , \4132 );
mnor \mul_7_15_g35422/U$1 ( \4512 , \4511 , \4464 );
mnor \mul_7_15_g35173/U$1 ( \4513 , \4510 , \4512 );
mnot \mul_7_15_g35172/U$1 ( \4514 , \4513 );
mnot \mul_7_15_g34778/U$3 ( \4515 , \4514 );
mnot \mul_7_15_g35606/U$3 ( \4516 , \4066 );
mnot \mul_7_15_g35606/U$4 ( \4517 , \4388 );
mor \mul_7_15_g35606/U$2 ( \4518 , \4516 , \4517 );
mnot \mul_7_15_g35947/U$1 ( \4519 , \4066 );
mnand \mul_7_15_g35884/U$1 ( \4520 , \4100 , \4519 );
mnand \mul_7_15_g35606/U$1 ( \4521 , \4518 , \4520 );
mnot \mul_7_15_g35068/U$3 ( \4522 , \4521 );
mnot \fopt36847/U$1 ( \4523 , \4193 );
mnot \mul_7_15_g35068/U$4 ( \4524 , \4523 );
mor \mul_7_15_g35068/U$2 ( \4525 , \4522 , \4524 );
mnand \mul_7_15_g35258/U$1 ( \4526 , \4393 , \4200 );
mnand \mul_7_15_g35068/U$1 ( \4527 , \4525 , \4526 );
mnot \mul_7_15_g34778/U$4 ( \4528 , \4527 );
mor \mul_7_15_g34778/U$2 ( \4529 , \4515 , \4528 );
mor \mul_7_15_g34880/U$2 ( \4530 , \4514 , \4527 );
mnot \mul_7_15_g35612/U$3 ( \4531 , \4051 );
mnot \mul_7_15_fopt36228/U$1 ( \4532 , \4458 );
mnot \mul_7_15_g35612/U$4 ( \4533 , \4532 );
mor \mul_7_15_g35612/U$2 ( \4534 , \4531 , \4533 );
mnot \mul_7_15_fopt36238/U$1 ( \4535 , \4436 );
mnot \mul_7_15_fopt36235/U$1 ( \4536 , \4535 );
mnand \mul_7_15_g35788/U$1 ( \4537 , \4536 , \4135 );
mnand \mul_7_15_g35612/U$1 ( \4538 , \4534 , \4537 );
mnot \mul_7_15_g35242/U$3 ( \4539 , \4538 );
mnot \mul_7_15_g35318/U$1 ( \4540 , \4450 );
mnot \mul_7_15_g35242/U$4 ( \4541 , \4540 );
mor \mul_7_15_g35242/U$2 ( \4542 , \4539 , \4541 );
mnot \mul_7_15_g35490/U$2 ( \4543 , \4532 );
mnand \mul_7_15_g35490/U$1 ( \4544 , \4543 , \4453 );
mnand \mul_7_15_g35242/U$1 ( \4545 , \4542 , \4544 );
mnand \mul_7_15_g34880/U$1 ( \4546 , \4530 , \4545 );
mnand \mul_7_15_g34778/U$1 ( \4547 , \4529 , \4546 );
mnand \mul_7_15_g34719/U$1 ( \4548 , \4503 , \4547 );
mnand \mul_7_15_g34738/U$1 ( \4549 , \4491 , \4502 );
mnand \mul_7_15_g34683/U$1 ( \4550 , \4548 , \4549 );
mxor \mul_7_15_g34569/U$1 ( \4551 , \4423 , \4473 );
mxor \mul_7_15_g34569/U$1_r1 ( \4552 , \4551 , \4484 );
mxor \mul_7_15_g34433/U$4 ( \4553 , \4550 , \4552 );
mxor \mul_7_15_g34808/U$1 ( \4554 , \4434 , \4459 );
mxor \mul_7_15_g34808/U$1_r1 ( \4555 , \4554 , \4470 );
mnot \mul_7_15_g36389/U$2 ( \4556 , \4555 );
mnot \mul_7_15_g35695/U$3 ( \4557 , \4096 );
mnot \mul_7_15_g35695/U$4 ( \4558 , \4163 );
mor \mul_7_15_g35695/U$2 ( \4559 , \4557 , \4558 );
mnand \mul_7_15_g35793/U$1 ( \4560 , \4170 , \4372 );
mnand \mul_7_15_g35695/U$1 ( \4561 , \4559 , \4560 );
mnot \mul_7_15_g35187/U$3 ( \4562 , \4561 );
mnot \mul_7_15_g35187/U$4 ( \4563 , \4159 );
mor \mul_7_15_g35187/U$2 ( \4564 , \4562 , \4563 );
mnand \mul_7_15_g35338/U$1 ( \4565 , \4150 , \4406 );
mnand \mul_7_15_g35187/U$1 ( \4566 , \4564 , \4565 );
mnot \mul_7_15_g35186/U$1 ( \4567 , \4566 );
mnand \mul_7_15_g35776/U$1 ( \4568 , \4102 , \4017 );
mnand \mul_7_15_g34992/U$1 ( \4569 , \4567 , \4568 );
mnot \mul_7_15_g35209/U$1 ( \4570 , \4502 );
mand \mul_7_15_g34851/U$2 ( \4571 , \4569 , \4570 );
mnor \mul_7_15_g34990/U$1 ( \4572 , \4567 , \4568 );
mnor \mul_7_15_g34851/U$1 ( \4573 , \4571 , \4572 );
mnand \mul_7_15_g36389/U$1 ( \4574 , \4556 , \4573 );
mnot \mul_7_15_g34534/U$3 ( \4575 , \4574 );
mxor \mul_7_15_g34633/U$1 ( \4576 , \4502 , \4547 );
mxnor \mul_7_15_g34633/U$1_r1 ( \4577 , \4576 , \4491 );
mnot \mul_7_15_g34587/U$1 ( \4578 , \4577 );
mnot \mul_7_15_g34534/U$4 ( \4579 , \4578 );
mor \mul_7_15_g34534/U$2 ( \4580 , \4575 , \4579 );
mnot \mul_7_15_g36384/U$2 ( \4581 , \4573 );
mnand \mul_7_15_g36384/U$1 ( \4582 , \4581 , \4555 );
mnand \mul_7_15_g34534/U$1 ( \4583 , \4580 , \4582 );
mand \mul_7_15_g34433/U$3 ( \4584 , \4553 , \4583 );
mand \mul_7_15_g34433/U$5 ( \4585 , \4550 , \4552 );
mor \mul_7_15_g34433/U$2 ( \4586 , \4584 , \4585 );
mnot \fopt36715/U$1 ( \4587 , \4586 );
mnand \mul_7_15_g34401/U$1 ( \4588 , \4489 , \4587 );
mbuf \mul_7_15_g34400/U$1 ( \4589 , \4588 );
mnot \mul_7_15_g36362/U$2 ( \4590 , \4589 );
mnot \mul_7_15_g34964/U$3 ( \4591 , \4513 );
mnot \mul_7_15_g34964/U$4 ( \4592 , \4527 );
mor \mul_7_15_g34964/U$2 ( \4593 , \4591 , \4592 );
mor \mul_7_15_g34964/U$5 ( \4594 , \4527 , \4513 );
mnand \mul_7_15_g34964/U$1 ( \4595 , \4593 , \4594 );
mxor \mul_7_15_g36417/U$1 ( \4596 , \4595 , \4545 );
mnot \mul_7_15_g35905/U$1 ( \4597 , \3516 );
mand \mul_7_15_g35539/U$2 ( \4598 , \2945 , \4597 );
mnot \mul_7_15_g35539/U$4 ( \4599 , \2945 );
mand \mul_7_15_g35539/U$3 ( \4600 , \4599 , \3516 );
mnor \mul_7_15_g35539/U$1 ( \4601 , \4598 , \4600 );
mbuf \mul_7_15_fopt36309/U$1 ( \4602 , \4601 );
mnot \mul_7_15_g35031/U$3 ( \4603 , \4602 );
mnot \mul_7_15_g35550/U$3 ( \4604 , \4442 );
mnot \mul_7_15_g35550/U$4 ( \4605 , \3516 );
mor \mul_7_15_g35550/U$2 ( \4606 , \4604 , \4605 );
mnand \mul_7_15_g35762/U$1 ( \4607 , \4597 , \3448 );
mnand \mul_7_15_g35550/U$1 ( \4608 , \4606 , \4607 );
mnand \mul_7_15_g35450/U$1 ( \4609 , \4608 , \4601 );
mnot \mul_7_15_g35449/U$1 ( \4610 , \4609 );
mbuf \mul_7_15_g35448/U$1 ( \4611 , \4610 );
mnot \mul_7_15_g35447/U$1 ( \4612 , \4611 );
mnot \mul_7_15_g35031/U$4 ( \4613 , \4612 );
mor \mul_7_15_g35031/U$2 ( \4614 , \4603 , \4613 );
mbuf \mul_7_15_g36149/U$1 ( \4615 , \3448 );
mbuf \mul_7_15_g36146/U$1 ( \4616 , \4615 );
mnand \mul_7_15_g35031/U$1 ( \4617 , \4614 , \4616 );
mnot \mul_7_15_g34906/U$3 ( \4618 , \4617 );
mnot \mul_7_15_g35218/U$3 ( \4619 , \4159 );
mnot \mul_7_15_g35687/U$3 ( \4620 , \4097 );
mnot \mul_7_15_g35687/U$4 ( \4621 , \4163 );
mor \mul_7_15_g35687/U$2 ( \4622 , \4620 , \4621 );
mnand \mul_7_15_g35825/U$1 ( \4623 , \4170 , \4254 );
mnand \mul_7_15_g35687/U$1 ( \4624 , \4622 , \4623 );
mnot \mul_7_15_g35218/U$4 ( \4625 , \4624 );
mor \mul_7_15_g35218/U$2 ( \4626 , \4619 , \4625 );
mnand \mul_7_15_g35377/U$1 ( \4627 , \4561 , \4150 );
mnand \mul_7_15_g35218/U$1 ( \4628 , \4626 , \4627 );
mnot \mul_7_15_g34906/U$4 ( \4629 , \4628 );
mor \mul_7_15_g34906/U$2 ( \4630 , \4618 , \4629 );
mor \mul_7_15_g34936/U$2 ( \4631 , \4628 , \4617 );
mbuf \mul_7_15_g35321/U$1 ( \4632 , \4449 );
mnot \mul_7_15_g35725/U$3 ( \4633 , \3997 );
mnot \mul_7_15_g35725/U$4 ( \4634 , \4535 );
mor \mul_7_15_g35725/U$2 ( \4635 , \4633 , \4634 );
mnand \mul_7_15_g35843/U$1 ( \4636 , \4536 , \4111 );
mnand \mul_7_15_g35725/U$1 ( \4637 , \4635 , \4636 );
mand \mul_7_15_g35083/U$2 ( \4638 , \4632 , \4637 );
mand \mul_7_15_g35083/U$3 ( \4639 , \4538 , \4453 );
mnor \mul_7_15_g35083/U$1 ( \4640 , \4638 , \4639 );
mnot \mul_7_15_g35082/U$1 ( \4641 , \4640 );
mnand \mul_7_15_g34936/U$1 ( \4642 , \4631 , \4641 );
mnand \mul_7_15_g34906/U$1 ( \4643 , \4630 , \4642 );
mxor \mul_7_15_g34596/U$4 ( \4644 , \4596 , \4643 );
mnot \mul_7_15_g35702/U$3 ( \4645 , \4095 );
mnot \mul_7_15_g35702/U$4 ( \4646 , \4134 );
mor \mul_7_15_g35702/U$2 ( \4647 , \4645 , \4646 );
mnand \mul_7_15_g35866/U$1 ( \4648 , \4106 , \4391 );
mnand \mul_7_15_g35702/U$1 ( \4649 , \4647 , \4648 );
mnot \mul_7_15_g35081/U$3 ( \4650 , \4649 );
mnot \mul_7_15_g35081/U$4 ( \4651 , \4302 );
mor \mul_7_15_g35081/U$2 ( \4652 , \4650 , \4651 );
mnot \mul_7_15_g36438/U$2 ( \4653 , \4507 );
mnot \mul_7_15_g35559/U$1 ( \4654 , \4511 );
mnand \mul_7_15_g36438/U$1 ( \4655 , \4653 , \4654 );
mnand \mul_7_15_g35081/U$1 ( \4656 , \4652 , \4655 );
mnot \mul_7_15_g35073/U$3 ( \4657 , \4395 );
mnot \mul_7_15_g35601/U$3 ( \4658 , \4017 );
mnot \mul_7_15_g35601/U$4 ( \4659 , \4101 );
mor \mul_7_15_g35601/U$2 ( \4660 , \4658 , \4659 );
mnot \mul_7_15_fopt36189/U$1 ( \4661 , \4346 );
mnot \mul_7_15_g36026/U$1 ( \4662 , \4017 );
mnand \mul_7_15_g36902/U$1 ( \4663 , \4661 , \4662 );
mnand \mul_7_15_g35601/U$1 ( \4664 , \4660 , \4663 );
mnot \mul_7_15_g35073/U$4 ( \4665 , \4664 );
mor \mul_7_15_g35073/U$2 ( \4666 , \4657 , \4665 );
mnand \mul_7_15_g35251/U$1 ( \4667 , \4521 , \4200 );
mnand \mul_7_15_g35073/U$1 ( \4668 , \4666 , \4667 );
mor \g37226/U$2 ( \4669 , \4656 , \4668 );
mnot \mul_7_15_g35663/U$3 ( \4670 , \4094 );
mnot \mul_7_15_g35663/U$4 ( \4671 , \4284 );
mor \mul_7_15_g35663/U$2 ( \4672 , \4670 , \4671 );
mnot \fopt36790/U$1 ( \4673 , \4332 );
mnand \mul_7_15_g35860/U$1 ( \4674 , \4673 , \4298 );
mnand \mul_7_15_g35663/U$1 ( \4675 , \4672 , \4674 );
mnot \mul_7_15_g35211/U$3 ( \4676 , \4675 );
mnot \mul_7_15_g35211/U$4 ( \4677 , \4430 );
mor \mul_7_15_g35211/U$2 ( \4678 , \4676 , \4677 );
mnand \mul_7_15_g35329/U$1 ( \4679 , \4497 , \4341 );
mnand \mul_7_15_g35211/U$1 ( \4680 , \4678 , \4679 );
mnand \g37226/U$1 ( \4681 , \4669 , \4680 );
mnot \fopt37227/U$1 ( \4682 , \4656 );
mnot \g37075/U$2 ( \4683 , \4682 );
mnand \g37075/U$1 ( \4684 , \4683 , \4668 );
mnand \g37225/U$1 ( \4685 , \4681 , \4684 );
mand \mul_7_15_g34596/U$3 ( \4686 , \4644 , \4685 );
mand \mul_7_15_g34596/U$5 ( \4687 , \4596 , \4643 );
mor \mul_7_15_g34596/U$2 ( \4688 , \4686 , \4687 );
mnot \mul_7_15_g34687/U$3 ( \4689 , \4573 );
mnot \mul_7_15_g34687/U$4 ( \4690 , \4555 );
mor \mul_7_15_g34687/U$2 ( \4691 , \4689 , \4690 );
mor \mul_7_15_g34687/U$5 ( \4692 , \4573 , \4555 );
mnand \mul_7_15_g34687/U$1 ( \4693 , \4691 , \4692 );
mnot \fopt36962/U$1 ( \4694 , \4693 );
mnot \mul_7_15_g34539/U$3 ( \4695 , \4694 );
mnot \mul_7_15_g34539/U$4 ( \4696 , \4578 );
mor \mul_7_15_g34539/U$2 ( \4697 , \4695 , \4696 );
mnand \mul_7_15_g34554/U$1 ( \4698 , \4577 , \4693 );
mnand \mul_7_15_g34539/U$1 ( \4699 , \4697 , \4698 );
mxor \mul_7_15_g34388/U$4 ( \4700 , \4688 , \4699 );
mxor \mul_7_15_g34856/U$1 ( \4701 , \4568 , \4566 );
mxnor \mul_7_15_g34856/U$1_r1 ( \4702 , \4701 , \4570 );
mnot \mul_7_15_g36383/U$2 ( \4703 , \4702 );
mnot \mul_7_15_g35647/U$3 ( \4704 , \4066 );
mnot \mul_7_15_g35647/U$4 ( \4705 , \4134 );
mor \mul_7_15_g35647/U$2 ( \4706 , \4704 , \4705 );
mnand \mul_7_15_g37187/U$1 ( \4707 , \4106 , \4519 );
mnand \mul_7_15_g35647/U$1 ( \4708 , \4706 , \4707 );
mnot \mul_7_15_g35107/U$3 ( \4709 , \4708 );
mnot \mul_7_15_g35451/U$1 ( \4710 , \4127 );
mnot \mul_7_15_g35107/U$4 ( \4711 , \4710 );
mor \mul_7_15_g35107/U$2 ( \4712 , \4709 , \4711 );
mnand \mul_7_15_g35373/U$1 ( \4713 , \4654 , \4649 );
mnand \mul_7_15_g35107/U$1 ( \4714 , \4712 , \4713 );
mnot \mul_7_15_g34785/U$3 ( \4715 , \4714 );
mnot \mul_7_15_g35670/U$3 ( \4716 , \4093 );
mnot \mul_7_15_g35670/U$4 ( \4717 , \4163 );
mor \mul_7_15_g35670/U$2 ( \4718 , \4716 , \4717 );
mnand \mul_7_15_g35839/U$1 ( \4719 , \4170 , \4349 );
mnand \mul_7_15_g35670/U$1 ( \4720 , \4718 , \4719 );
mnot \mul_7_15_g35124/U$3 ( \4721 , \4720 );
mnot \mul_7_15_g35124/U$4 ( \4722 , \4159 );
mor \mul_7_15_g35124/U$2 ( \4723 , \4721 , \4722 );
mnand \mul_7_15_g35351/U$1 ( \4724 , \4624 , \4317 );
mnand \mul_7_15_g35124/U$1 ( \4725 , \4723 , \4724 );
mnot \mul_7_15_g34785/U$4 ( \4726 , \4725 );
mor \mul_7_15_g34785/U$2 ( \4727 , \4715 , \4726 );
mor \mul_7_15_g34870/U$2 ( \4728 , \4714 , \4725 );
mbuf \mul_7_15_fopt36241/U$1 ( \4729 , \4436 );
mand \mul_7_15_g35641/U$2 ( \4730 , \4198 , \4729 );
mnot \mul_7_15_g35641/U$4 ( \4731 , \4198 );
mbuf \mul_7_15_fopt36224/U$1 ( \4732 , \4457 );
mand \mul_7_15_g35641/U$3 ( \4733 , \4731 , \4732 );
mnor \mul_7_15_g35641/U$1 ( \4734 , \4730 , \4733 );
mnot \mul_7_15_g35103/U$3 ( \4735 , \4734 );
mnot \mul_7_15_g35103/U$4 ( \4736 , \4540 );
mor \mul_7_15_g35103/U$2 ( \4737 , \4735 , \4736 );
mnand \mul_7_15_g35353/U$1 ( \4738 , \4637 , \4453 );
mnand \mul_7_15_g35103/U$1 ( \4739 , \4737 , \4738 );
mnand \mul_7_15_g34870/U$1 ( \4740 , \4728 , \4739 );
mnand \mul_7_15_g34785/U$1 ( \4741 , \4727 , \4740 );
mand \mul_7_15_g35781/U$1 ( \4742 , \4102 , \4021 );
mnot \mul_7_15_g36425/U$2 ( \4743 , \4742 );
mnot \mul_7_15_g35613/U$3 ( \4744 , \4051 );
mbuf \mul_7_15_g36135/U$1 ( \4745 , \3448 );
mnot \mul_7_15_g36132/U$1 ( \4746 , \4745 );
mnot \mul_7_15_g35613/U$4 ( \4747 , \4746 );
mor \mul_7_15_g35613/U$2 ( \4748 , \4744 , \4747 );
mnand \mul_7_15_g35789/U$1 ( \4749 , \4745 , \4135 );
mnand \mul_7_15_g35613/U$1 ( \4750 , \4748 , \4749 );
mnot \mul_7_15_g35239/U$3 ( \4751 , \4750 );
mnot \mul_7_15_g35239/U$4 ( \4752 , \4611 );
mor \mul_7_15_g35239/U$2 ( \4753 , \4751 , \4752 );
mnot \mul_7_15_fopt36307/U$1 ( \4754 , \4602 );
mnand \mul_7_15_g35489/U$1 ( \4755 , \4754 , \4616 );
mnand \mul_7_15_g35239/U$1 ( \4756 , \4753 , \4755 );
mnot \mul_7_15_g35238/U$1 ( \4757 , \4756 );
mnand \mul_7_15_g36425/U$1 ( \4758 , \4743 , \4757 );
mand \mul_7_15_g34686/U$2 ( \4759 , \4741 , \4758 );
mand \mul_7_15_g34920/U$2 ( \4760 , \4742 , \4756 );
mnor \mul_7_15_g34686/U$1 ( \4761 , \4759 , \4760 );
mnand \mul_7_15_g36383/U$1 ( \4762 , \4703 , \4761 );
mnot \mul_7_15_g34509/U$3 ( \4763 , \4762 );
mand \g37074/U$2 ( \4764 , \4680 , \4656 );
mnot \g37074/U$4 ( \4765 , \4680 );
mand \g37074/U$3 ( \4766 , \4765 , \4682 );
mnor \g37074/U$1 ( \4767 , \4764 , \4766 );
mnot \mul_7_15_g37228/U$1 ( \4768 , \4668 );
mand \mul_7_15_g34893/U$2 ( \4769 , \4767 , \4768 );
mnot \mul_7_15_g34893/U$4 ( \4770 , \4767 );
mand \mul_7_15_g34893/U$3 ( \4771 , \4770 , \4668 );
mnor \mul_7_15_g34893/U$1 ( \4772 , \4769 , \4771 );
mnot \mul_7_15_fopt36310/U$1 ( \4773 , \4772 );
mnot \g37146/U$3 ( \4774 , \4773 );
mand \mul_7_15_g36352/U$1 ( \4775 , \4100 , \4026 );
mnot \mul_7_15_g34928/U$3 ( \4776 , \4775 );
mnot \mul_7_15_g35598/U$3 ( \4777 , \4021 );
mnot \mul_7_15_g35598/U$4 ( \4778 , \4101 );
mor \mul_7_15_g35598/U$2 ( \4779 , \4777 , \4778 );
mnot \mul_7_15_g36024/U$1 ( \4780 , \4021 );
mnand \mul_7_15_g35856/U$1 ( \4781 , \4100 , \4780 );
mnand \mul_7_15_g35598/U$1 ( \4782 , \4779 , \4781 );
mnot \mul_7_15_g35058/U$3 ( \4783 , \4782 );
mnot \mul_7_15_g35058/U$4 ( \4784 , \4395 );
mor \mul_7_15_g35058/U$2 ( \4785 , \4783 , \4784 );
mnand \mul_7_15_g35253/U$1 ( \4786 , \4664 , \4200 );
mnand \mul_7_15_g35058/U$1 ( \4787 , \4785 , \4786 );
mnot \mul_7_15_g34928/U$4 ( \4788 , \4787 );
mor \mul_7_15_g34928/U$2 ( \4789 , \4776 , \4788 );
mor \mul_7_15_g34941/U$2 ( \4790 , \4787 , \4775 );
mnot \mul_7_15_g35631/U$3 ( \4791 , \4096 );
mnot \mul_7_15_g35631/U$4 ( \4792 , \4284 );
mor \mul_7_15_g35631/U$2 ( \4793 , \4791 , \4792 );
mnand \mul_7_15_g35792/U$1 ( \4794 , \4283 , \4372 );
mnand \mul_7_15_g35631/U$1 ( \4795 , \4793 , \4794 );
mnot \mul_7_15_g35091/U$3 ( \4796 , \4795 );
mnot \fopt36696/U$1 ( \4797 , \4278 );
mnot \mul_7_15_g35091/U$4 ( \4798 , \4797 );
mor \mul_7_15_g35091/U$2 ( \4799 , \4796 , \4798 );
mnot \mul_7_15_g35575/U$1 ( \4800 , \4265 );
mnand \mul_7_15_g35348/U$1 ( \4801 , \4675 , \4800 );
mnand \mul_7_15_g35091/U$1 ( \4802 , \4799 , \4801 );
mnand \mul_7_15_g34941/U$1 ( \4803 , \4790 , \4802 );
mnand \mul_7_15_g34928/U$1 ( \4804 , \4789 , \4803 );
mnot \g37146/U$4 ( \4805 , \4804 );
mor \g37146/U$2 ( \4806 , \4774 , \4805 );
mnot \mul_7_15_g34845/U$1 ( \4807 , \4804 );
mnot \g37147/U$3 ( \4808 , \4807 );
mnot \g37147/U$4 ( \4809 , \4772 );
mor \g37147/U$2 ( \4810 , \4808 , \4809 );
mxor \g36562/U$1 ( \4811 , \4617 , \4640 );
mxnor \g36562/U$1_r1 ( \4812 , \4811 , \4628 );
mnand \g37147/U$1 ( \4813 , \4810 , \4812 );
mnand \g37146/U$1 ( \4814 , \4806 , \4813 );
mnot \mul_7_15_g34509/U$4 ( \4815 , \4814 );
mor \mul_7_15_g34509/U$2 ( \4816 , \4763 , \4815 );
mnot \mul_7_15_g36378/U$2 ( \4817 , \4761 );
mnand \mul_7_15_g36378/U$1 ( \4818 , \4817 , \4702 );
mnand \mul_7_15_g34509/U$1 ( \4819 , \4816 , \4818 );
mand \mul_7_15_g34388/U$3 ( \4820 , \4700 , \4819 );
mand \mul_7_15_g34388/U$5 ( \4821 , \4688 , \4699 );
mor \mul_7_15_g34388/U$2 ( \4822 , \4820 , \4821 );
mxor \mul_7_15_g34433/U$1 ( \4823 , \4550 , \4552 );
mxor \mul_7_15_g34433/U$1_r1 ( \4824 , \4823 , \4583 );
mnor \mul_7_15_g34354/U$1 ( \4825 , \4822 , \4824 );
mnot \mul_7_15_g34319/U$2 ( \4826 , \4825 );
mxor \mul_7_15_g34388/U$1 ( \4827 , \4688 , \4699 );
mxor \mul_7_15_g34388/U$1_r1 ( \4828 , \4827 , \4819 );
mnot \mul_7_15_g34583/U$3 ( \4829 , \4761 );
mnot \mul_7_15_g34583/U$4 ( \4830 , \4702 );
mor \mul_7_15_g34583/U$2 ( \4831 , \4829 , \4830 );
mor \mul_7_15_g34583/U$5 ( \4832 , \4761 , \4702 );
mnand \mul_7_15_g34583/U$1 ( \4833 , \4831 , \4832 );
mxor \g37092/U$1 ( \4834 , \4814 , \4833 );
mnot \g37091/U$3 ( \4835 , \4834 );
mxor \mul_7_15_g34596/U$1 ( \4836 , \4596 , \4643 );
mxor \mul_7_15_g34596/U$1_r1 ( \4837 , \4836 , \4685 );
mbuf \mul_7_15_g34595/U$1 ( \4838 , \4837 );
mnot \g37091/U$4 ( \4839 , \4838 );
mor \g37091/U$2 ( \4840 , \4835 , \4839 );
mor \mul_7_15_g34407/U$2 ( \4841 , \4838 , \4834 );
mxor \mul_7_15_g34920/U$1 ( \4842 , \4742 , \4756 );
mand \mul_7_15_g34688/U$2 ( \4843 , \4741 , \4842 );
mnot \mul_7_15_g34688/U$4 ( \4844 , \4741 );
mnot \mul_7_15_g34919/U$1 ( \4845 , \4842 );
mand \mul_7_15_g34688/U$3 ( \4846 , \4844 , \4845 );
mnor \mul_7_15_g34688/U$1 ( \4847 , \4843 , \4846 );
mbuf \mul_7_15_g34673/U$1 ( \4848 , \4847 );
mnot \mul_7_15_g34447/U$3 ( \4849 , \4848 );
mnot \mul_7_15_g34579/U$3 ( \4850 , \4757 );
mbuf \mul_7_15_g35951/U$1 ( \4851 , \3016 );
mnot \mul_7_15_g35552/U$3 ( \4852 , \4851 );
mnot \mul_7_15_g35973/U$1 ( \4853 , \2945 );
mnot \mul_7_15_g35552/U$4 ( \4854 , \4853 );
mor \mul_7_15_g35552/U$2 ( \4855 , \4852 , \4854 );
mnot \mul_7_15_g35948/U$1 ( \4856 , \4851 );
mnand \mul_7_15_g35765/U$1 ( \4857 , \4856 , \2945 );
mnand \mul_7_15_g35552/U$1 ( \4858 , \4855 , \4857 );
mbuf \mul_7_15_g35551/U$1 ( \4859 , \4858 );
mnot \mul_7_15_g35269/U$3 ( \4860 , \4859 );
mxnor \g36556/U$1 ( \4861 , \3016 , \3070 );
mbuf \mul_7_15_fopt36164/U$1 ( \4862 , \4861 );
mnot \mul_7_15_fopt36155/U$1 ( \4863 , \4862 );
mnot \mul_7_15_g35269/U$4 ( \4864 , \4863 );
mand \mul_7_15_g35269/U$2 ( \4865 , \4860 , \4864 );
mbuf \mul_7_15_g35969/U$1 ( \4866 , \4853 );
mnot \mul_7_15_g35967/U$1 ( \4867 , \4866 );
mbuf \mul_7_15_g35966/U$1 ( \4868 , \4867 );
mnot \mul_7_15_g35963/U$1 ( \4869 , \4868 );
mnor \mul_7_15_g35269/U$1 ( \4870 , \4865 , \4869 );
mnot \mul_7_15_g35268/U$1 ( \4871 , \4870 );
mnot \mul_7_15_g34784/U$3 ( \4872 , \4871 );
mnot \mul_7_15_g35121/U$3 ( \4873 , \4610 );
mnot \mul_7_15_g35645/U$3 ( \4874 , \3997 );
mnot \mul_7_15_g35645/U$4 ( \4875 , \4746 );
mor \mul_7_15_g35645/U$2 ( \4876 , \4874 , \4875 );
mnand \mul_7_15_g35832/U$1 ( \4877 , \4745 , \4111 );
mnand \mul_7_15_g35645/U$1 ( \4878 , \4876 , \4877 );
mnot \mul_7_15_g35121/U$4 ( \4879 , \4878 );
mor \mul_7_15_g35121/U$2 ( \4880 , \4873 , \4879 );
mnot \mul_7_15_fopt36300/U$1 ( \4881 , \4602 );
mnand \mul_7_15_g35440/U$1 ( \4882 , \4881 , \4750 );
mnand \mul_7_15_g35121/U$1 ( \4883 , \4880 , \4882 );
mnot \mul_7_15_g34784/U$4 ( \4884 , \4883 );
mor \mul_7_15_g34784/U$2 ( \4885 , \4872 , \4884 );
mor \mul_7_15_g34876/U$2 ( \4886 , \4871 , \4883 );
mnot \mul_7_15_g35662/U$3 ( \4887 , \4097 );
mnot \mul_7_15_g35662/U$4 ( \4888 , \4493 );
mor \mul_7_15_g35662/U$2 ( \4889 , \4887 , \4888 );
mnand \mul_7_15_g35799/U$1 ( \4890 , \4285 , \4254 );
mnand \mul_7_15_g35662/U$1 ( \4891 , \4889 , \4890 );
mnot \mul_7_15_g35123/U$3 ( \4892 , \4891 );
mnot \mul_7_15_g35123/U$4 ( \4893 , \4430 );
mor \mul_7_15_g35123/U$2 ( \4894 , \4892 , \4893 );
mnand \mul_7_15_g35367/U$1 ( \4895 , \4341 , \4795 );
mnand \mul_7_15_g35123/U$1 ( \4896 , \4894 , \4895 );
mnand \mul_7_15_g34876/U$1 ( \4897 , \4886 , \4896 );
mnand \mul_7_15_g34784/U$1 ( \4898 , \4885 , \4897 );
mnot \mul_7_15_g34579/U$4 ( \4899 , \4898 );
mor \mul_7_15_g34579/U$2 ( \4900 , \4850 , \4899 );
mor \mul_7_15_g34619/U$2 ( \4901 , \4757 , \4898 );
mand \mul_7_15_g35777/U$1 ( \4902 , \4102 , \4072 );
mnot \mul_7_15_g34794/U$3 ( \4903 , \4902 );
mnot \mul_7_15_g35665/U$3 ( \4904 , \4095 );
mnot \mul_7_15_g35665/U$4 ( \4905 , \4163 );
mor \mul_7_15_g35665/U$2 ( \4906 , \4904 , \4905 );
mnand \mul_7_15_g35885/U$1 ( \4907 , \4164 , \4391 );
mnand \mul_7_15_g35665/U$1 ( \4908 , \4906 , \4907 );
mnot \mul_7_15_g35126/U$3 ( \4909 , \4908 );
mnot \mul_7_15_g35126/U$4 ( \4910 , \4159 );
mor \mul_7_15_g35126/U$2 ( \4911 , \4909 , \4910 );
mnand \mul_7_15_g35371/U$1 ( \4912 , \4150 , \4720 );
mnand \mul_7_15_g35126/U$1 ( \4913 , \4911 , \4912 );
mnot \mul_7_15_g34794/U$4 ( \4914 , \4913 );
mor \mul_7_15_g34794/U$2 ( \4915 , \4903 , \4914 );
mor \mul_7_15_g34877/U$2 ( \4916 , \4913 , \4902 );
mnot \mul_7_15_fopt36223/U$1 ( \4917 , \4732 );
mand \mul_7_15_g35666/U$2 ( \4918 , \4094 , \4917 );
mnot \mul_7_15_g35666/U$4 ( \4919 , \4094 );
mand \mul_7_15_g35666/U$3 ( \4920 , \4919 , \4535 );
mnor \mul_7_15_g35666/U$1 ( \4921 , \4918 , \4920 );
mnot \mul_7_15_g35131/U$3 ( \4922 , \4921 );
mnot \mul_7_15_g35131/U$4 ( \4923 , \4632 );
mor \mul_7_15_g35131/U$2 ( \4924 , \4922 , \4923 );
mnand \mul_7_15_g35366/U$1 ( \4925 , \4453 , \4734 );
mnand \mul_7_15_g35131/U$1 ( \4926 , \4924 , \4925 );
mnand \mul_7_15_g34877/U$1 ( \4927 , \4916 , \4926 );
mnand \mul_7_15_g34794/U$1 ( \4928 , \4915 , \4927 );
mnand \mul_7_15_g34619/U$1 ( \4929 , \4901 , \4928 );
mnand \mul_7_15_g34579/U$1 ( \4930 , \4900 , \4929 );
mnot \mul_7_15_g34447/U$4 ( \4931 , \4930 );
mor \mul_7_15_g34447/U$2 ( \4932 , \4849 , \4931 );
mor \mul_7_15_g34468/U$2 ( \4933 , \4848 , \4930 );
mbuf \mul_7_15_g35989/U$1 ( \4934 , \2945 );
mnot \mul_7_15_g35988/U$1 ( \4935 , \4934 );
mnot \mul_7_15_g35986/U$1 ( \4936 , \4935 );
mand \mul_7_15_g35611/U$2 ( \4937 , \4051 , \4936 );
mnot \mul_7_15_g35611/U$4 ( \4938 , \4051 );
mnot \mul_7_15_g35982/U$1 ( \4939 , \4934 );
mand \mul_7_15_g35611/U$3 ( \4940 , \4938 , \4939 );
mnor \mul_7_15_g35611/U$1 ( \4941 , \4937 , \4940 );
mnot \mul_7_15_g35233/U$3 ( \4942 , \4941 );
mnand \mul_7_15_g35471/U$1 ( \4943 , \4858 , \4862 );
mnot \mul_7_15_g35470/U$1 ( \4944 , \4943 );
mbuf \mul_7_15_g35469/U$1 ( \4945 , \4944 );
mnot \mul_7_15_g35233/U$4 ( \4946 , \4945 );
mor \mul_7_15_g35233/U$2 ( \4947 , \4942 , \4946 );
mnot \mul_7_15_fopt36157/U$1 ( \4948 , \4862 );
mnot \mul_7_15_g35981/U$1 ( \4949 , \4939 );
mnand \mul_7_15_g35486/U$1 ( \4950 , \4948 , \4949 );
mnand \mul_7_15_g35233/U$1 ( \4951 , \4947 , \4950 );
mnot \mul_7_15_g34916/U$3 ( \4952 , \4951 );
mnot \mul_7_15_g35640/U$3 ( \4953 , \4017 );
mnot \mul_7_15_g35640/U$4 ( \4954 , \4134 );
mor \mul_7_15_g35640/U$2 ( \4955 , \4953 , \4954 );
mnand \mul_7_15_g36693/U$1 ( \4956 , \4106 , \4662 );
mnand \mul_7_15_g35640/U$1 ( \4957 , \4955 , \4956 );
mnot \mul_7_15_g35140/U$3 ( \4958 , \4957 );
mnot \mul_7_15_g35140/U$4 ( \4959 , \4302 );
mor \mul_7_15_g35140/U$2 ( \4960 , \4958 , \4959 );
mnand \mul_7_15_g35444/U$1 ( \4961 , \4654 , \4708 );
mnand \mul_7_15_g35140/U$1 ( \4962 , \4960 , \4961 );
mnot \mul_7_15_g34916/U$4 ( \4963 , \4962 );
mor \mul_7_15_g34916/U$2 ( \4964 , \4952 , \4963 );
mor \mul_7_15_g34940/U$2 ( \4965 , \4951 , \4962 );
mnot \mul_7_15_g35607/U$3 ( \4966 , \4026 );
mnot \mul_7_15_g35607/U$4 ( \4967 , \4250 );
mor \mul_7_15_g35607/U$2 ( \4968 , \4966 , \4967 );
mnot \mul_7_15_g36027/U$1 ( \4969 , \4026 );
mnand \mul_7_15_g35824/U$1 ( \4970 , \4661 , \4969 );
mnand \mul_7_15_g35607/U$1 ( \4971 , \4968 , \4970 );
mnot \mul_7_15_g35062/U$3 ( \4972 , \4971 );
mnot \mul_7_15_g35062/U$4 ( \4973 , \4395 );
mor \mul_7_15_g35062/U$2 ( \4974 , \4972 , \4973 );
mnand \mul_7_15_g35260/U$1 ( \4975 , \4782 , \4200 );
mnand \mul_7_15_g35062/U$1 ( \4976 , \4974 , \4975 );
mnand \mul_7_15_g34940/U$1 ( \4977 , \4965 , \4976 );
mnand \mul_7_15_g34916/U$1 ( \4978 , \4964 , \4977 );
mnot \fopt36907/U$1 ( \4979 , \4978 );
mnot \mul_7_15_g34653/U$3 ( \4980 , \4979 );
mxor \mul_7_15_g34902/U$1 ( \4981 , \4775 , \4802 );
mxnor \mul_7_15_g34902/U$1_r1 ( \4982 , \4981 , \4787 );
mnot \mul_7_15_g34653/U$4 ( \4983 , \4982 );
mor \mul_7_15_g34653/U$2 ( \4984 , \4980 , \4983 );
mnot \mul_7_15_g34970/U$3 ( \4985 , \4725 );
mnot \mul_7_15_g35106/U$1 ( \4986 , \4714 );
mnot \mul_7_15_g34970/U$4 ( \4987 , \4986 );
mor \mul_7_15_g34970/U$2 ( \4988 , \4985 , \4987 );
mnot \mul_7_15_g34984/U$2 ( \4989 , \4725 );
mnand \mul_7_15_g34984/U$1 ( \4990 , \4989 , \4714 );
mnand \mul_7_15_g34970/U$1 ( \4991 , \4988 , \4990 );
mand \mul_7_15_g34858/U$2 ( \4992 , \4991 , \4739 );
mnot \mul_7_15_g34858/U$4 ( \4993 , \4991 );
mnot \fopt36857/U$1 ( \4994 , \4739 );
mand \mul_7_15_g34858/U$3 ( \4995 , \4993 , \4994 );
mnor \mul_7_15_g34858/U$1 ( \4996 , \4992 , \4995 );
mnand \mul_7_15_g34653/U$1 ( \4997 , \4984 , \4996 );
mor \mul_7_15_g36390/U$1 ( \4998 , \4982 , \4979 );
mnand \mul_7_15_g34628/U$1 ( \4999 , \4997 , \4998 );
mnand \mul_7_15_g34468/U$1 ( \5000 , \4933 , \4999 );
mnand \mul_7_15_g34447/U$1 ( \5001 , \4932 , \5000 );
mnand \mul_7_15_g34407/U$1 ( \5002 , \4841 , \5001 );
mnand \g37091/U$1 ( \5003 , \4840 , \5002 );
mor \mul_7_15_g36359/U$1 ( \5004 , \4828 , \5003 );
mnand \mul_7_15_g34319/U$1 ( \5005 , \4826 , \5004 );
mnor \mul_7_15_g36362/U$1 ( \5006 , \4590 , \5005 );
mxor \mul_7_15_g34452/U$4 ( \5007 , \4418 , \4420 );
mand \mul_7_15_g34452/U$3 ( \5008 , \5007 , \4487 );
mand \mul_7_15_g34452/U$5 ( \5009 , \4418 , \4420 );
mor \mul_7_15_g34452/U$2 ( \5010 , \5008 , \5009 );
mxor \mul_7_15_g36835/U$1 ( \5011 , \4322 , \4325 );
mxor \mul_7_15_g36835/U$1_r1 ( \5012 , \5011 , \4365 );
mor \mul_7_15_g34427/U$1 ( \5013 , \5010 , \5012 );
mnand \mul_7_15_g34267/U$1 ( \5014 , \5006 , \5013 );
mnor \mul_7_15_g36367/U$1 ( \5015 , \4371 , \5014 );
mor \g37270/U$2 ( \5016 , \4230 , \4166 );
mnand \g37270/U$1 ( \5017 , \5016 , \4292 );
mnand \mul_7_15_g34617/U$1 ( \5018 , \4166 , \4230 );
mnand \mul_7_15_g34510/U$1 ( \5019 , \5017 , \5018 );
mxor \mul_7_15_g34814/U$4 ( \5020 , \4103 , \4141 );
mand \mul_7_15_g34814/U$3 ( \5021 , \5020 , \4165 );
mand \mul_7_15_g34814/U$5 ( \5022 , \4103 , \4141 );
mor \mul_7_15_g34814/U$2 ( \5023 , \5021 , \5022 );
mand \mul_7_15_g35511/U$2 ( \5024 , \4094 , \4100 );
mnand \mul_7_15_g35248/U$1 ( \5025 , \4129 , \4139 );
mnand \mul_7_15_g35491/U$1 ( \5026 , \4133 , \4106 );
mand \mul_7_15_g35235/U$1 ( \5027 , \5025 , \5026 );
mxor \mul_7_15_g34823/U$1 ( \5028 , \5024 , \5027 );
mnot \fopt36852/U$1 ( \5029 , \4195 );
mnot \mul_7_15_g35515/U$1 ( \5030 , \4199 );
mor \mul_7_15_g35063/U$2 ( \5031 , \5029 , \5030 );
mand \g36923/U$2 ( \5032 , \4102 , \4111 );
mnot \g36923/U$4 ( \5033 , \4102 );
mand \g36923/U$3 ( \5034 , \5033 , \3997 );
mnor \g36923/U$1 ( \5035 , \5032 , \5034 );
mor \mul_7_15_g35063/U$3 ( \5036 , \5035 , \4192 );
mnand \mul_7_15_g35063/U$1 ( \5037 , \5031 , \5036 );
mxor \mul_7_15_g34823/U$1_r1 ( \5038 , \5028 , \5037 );
mxor \mul_7_15_g34565/U$1 ( \5039 , \5023 , \5038 );
mxor \mul_7_15_g34670/U$4 ( \5040 , \4177 , \4202 );
mand \mul_7_15_g34670/U$3 ( \5041 , \5040 , \4229 );
mand \mul_7_15_g34670/U$5 ( \5042 , \4177 , \4202 );
mor \mul_7_15_g34670/U$2 ( \5043 , \5041 , \5042 );
mxor \mul_7_15_g34565/U$1_r1 ( \5044 , \5039 , \5043 );
mor \mul_7_15_g36371/U$1 ( \5045 , \5019 , \5044 );
mnand \mul_7_15_g34231/U$1 ( \5046 , \5015 , \5045 );
mxor \mul_7_15_g34565/U$4 ( \5047 , \5023 , \5038 );
mand \mul_7_15_g34565/U$3 ( \5048 , \5047 , \5043 );
mand \mul_7_15_g34565/U$5 ( \5049 , \5023 , \5038 );
mor \mul_7_15_g34565/U$2 ( \5050 , \5048 , \5049 );
mnot \mul_7_15_g35234/U$1 ( \5051 , \5027 );
mxor \mul_7_15_g34823/U$4 ( \5052 , \5024 , \5027 );
mand \mul_7_15_g34823/U$3 ( \5053 , \5052 , \5037 );
mand \mul_7_15_g34823/U$5 ( \5054 , \5024 , \5027 );
mor \mul_7_15_g34823/U$2 ( \5055 , \5053 , \5054 );
mxor \mul_7_15_g34599/U$1 ( \5056 , \5051 , \5055 );
mand \mul_7_15_g35516/U$2 ( \5057 , \4198 , \4102 );
mor \mul_7_15_g36421/U$2 ( \5058 , \4133 , \4302 );
mnand \mul_7_15_g36421/U$1 ( \5059 , \5058 , \4106 );
mxor \mul_7_15_g34832/U$1 ( \5060 , \5057 , \5059 );
mor \mul_7_15_g35055/U$2 ( \5061 , \5029 , \5035 );
mand \mul_7_15_g35597/U$2 ( \5062 , \4101 , \4051 );
mand \mul_7_15_g35597/U$3 ( \5063 , \4102 , \4135 );
mnor \mul_7_15_g35597/U$1 ( \5064 , \5062 , \5063 );
mor \mul_7_15_g35055/U$3 ( \5065 , \5064 , \4192 );
mnand \mul_7_15_g35055/U$1 ( \5066 , \5061 , \5065 );
mxor \mul_7_15_g34832/U$1_r1 ( \5067 , \5060 , \5066 );
mxor \mul_7_15_g34599/U$1_r1 ( \5068 , \5056 , \5067 );
mnor \mul_7_15_g34522/U$1 ( \5069 , \5050 , \5068 );
mnor \mul_7_15_g34215/U$1 ( \5070 , \5046 , \5069 );
mnot \mul_7_15_g34187/U$3 ( \5071 , \5070 );
mxor \mul_7_15_g36408/U$1 ( \5072 , \4962 , \4976 );
mbuf \mul_7_15_g35231/U$1 ( \5073 , \4951 );
mnot \mul_7_15_g35230/U$1 ( \5074 , \5073 );
mand \mul_7_15_g34899/U$2 ( \5075 , \5072 , \5074 );
mnot \mul_7_15_g34899/U$4 ( \5076 , \5072 );
mand \mul_7_15_g34899/U$3 ( \5077 , \5076 , \5073 );
mnor \mul_7_15_g34899/U$1 ( \5078 , \5075 , \5077 );
mnot \mul_7_15_fopt36166/U$1 ( \5079 , \5078 );
mnot \mul_7_15_fopt36165/U$1 ( \5080 , \5079 );
mxor \mul_7_15_g36424/U$1 ( \5081 , \4913 , \4902 );
mbuf \fopt36705/U$1 ( \5082 , \4926 );
mxnor \mul_7_15_g36406/U$1 ( \5083 , \5081 , \5082 );
mnand \mul_7_15_g36439/U$1 ( \5084 , \5080 , \5083 );
mnot \mul_7_15_g34800/U$3 ( \5085 , \5074 );
mnot \mul_7_15_g35602/U$3 ( \5086 , \4072 );
mnot \mul_7_15_g35602/U$4 ( \5087 , \4250 );
mor \mul_7_15_g35602/U$2 ( \5088 , \5086 , \5087 );
mnot \mul_7_15_g35912/U$1 ( \5089 , \4072 );
mnand \mul_7_15_g35887/U$1 ( \5090 , \4661 , \5089 );
mnand \mul_7_15_g35602/U$1 ( \5091 , \5088 , \5090 );
mnot \mul_7_15_g35070/U$3 ( \5092 , \5091 );
mnot \mul_7_15_g35070/U$4 ( \5093 , \4395 );
mor \mul_7_15_g35070/U$2 ( \5094 , \5092 , \5093 );
mnand \mul_7_15_g35261/U$1 ( \5095 , \4971 , \4200 );
mnand \mul_7_15_g35070/U$1 ( \5096 , \5094 , \5095 );
mnot \mul_7_15_g34800/U$4 ( \5097 , \5096 );
mor \mul_7_15_g34800/U$2 ( \5098 , \5085 , \5097 );
mnot \mul_7_15_g34881/U$3 ( \5099 , \4951 );
mnot \mul_7_15_g35069/U$1 ( \5100 , \5096 );
mnot \mul_7_15_g34881/U$4 ( \5101 , \5100 );
mor \mul_7_15_g34881/U$2 ( \5102 , \5099 , \5101 );
mnot \mul_7_15_g35700/U$3 ( \5103 , \3997 );
mnot \mul_7_15_g35700/U$4 ( \5104 , \4939 );
mor \mul_7_15_g35700/U$2 ( \5105 , \5103 , \5104 );
mnand \mul_7_15_g35847/U$1 ( \5106 , \4867 , \4111 );
mnand \mul_7_15_g35700/U$1 ( \5107 , \5105 , \5106 );
mand \g37141/U$2 ( \5108 , \4945 , \5107 );
mand \g37141/U$3 ( \5109 , \4863 , \4941 );
mnor \g37141/U$1 ( \5110 , \5108 , \5109 );
mnot \mul_7_15_g35620/U$3 ( \5111 , \4097 );
mnot \mul_7_15_fopt36240/U$1 ( \5112 , \4729 );
mnot \mul_7_15_g35620/U$4 ( \5113 , \5112 );
mor \mul_7_15_g35620/U$2 ( \5114 , \5111 , \5113 );
mnand \mul_7_15_g35810/U$1 ( \5115 , \4458 , \4254 );
mnand \mul_7_15_g35620/U$1 ( \5116 , \5114 , \5115 );
mand \mul_7_15_g35194/U$2 ( \5117 , \5116 , \4632 );
mnot \mul_7_15_g35716/U$3 ( \5118 , \4096 );
mnot \mul_7_15_g35716/U$4 ( \5119 , \4535 );
mor \mul_7_15_g35716/U$2 ( \5120 , \5118 , \5119 );
mnand \mul_7_15_g35883/U$1 ( \5121 , \4536 , \4372 );
mnand \mul_7_15_g35716/U$1 ( \5122 , \5120 , \5121 );
mand \mul_7_15_g35194/U$3 ( \5123 , \5122 , \4453 );
mnor \mul_7_15_g35194/U$1 ( \5124 , \5117 , \5123 );
mnand \mul_7_15_g34988/U$1 ( \5125 , \5110 , \5124 );
mnand \mul_7_15_g34881/U$1 ( \5126 , \5102 , \5125 );
mnand \mul_7_15_g34800/U$1 ( \5127 , \5098 , \5126 );
mand \mul_7_15_g34656/U$2 ( \5128 , \5084 , \5127 );
mnor \mul_7_15_g34706/U$1 ( \5129 , \5080 , \5083 );
mnor \mul_7_15_g34656/U$1 ( \5130 , \5128 , \5129 );
mxor \mul_7_15_g34584/U$1 ( \5131 , \4757 , \4898 );
mxnor \mul_7_15_g34584/U$1_r1 ( \5132 , \5131 , \4928 );
mnot \mul_7_15_fopt36193/U$1 ( \5133 , \4250 );
mnand \mul_7_15_g35779/U$1 ( \5134 , \5133 , \4076 );
mnot \mul_7_15_g35778/U$1 ( \5135 , \5134 );
mnot \mul_7_15_g34795/U$3 ( \5136 , \5135 );
mnot \mul_7_15_g35703/U$3 ( \5137 , \4198 );
mnot \mul_7_15_g36143/U$1 ( \5138 , \4615 );
mnot \mul_7_15_g35703/U$4 ( \5139 , \5138 );
mor \mul_7_15_g35703/U$2 ( \5140 , \5137 , \5139 );
mnand \mul_7_15_g36927/U$1 ( \5141 , \4616 , \4209 );
mnand \mul_7_15_g35703/U$1 ( \5142 , \5140 , \5141 );
mnot \mul_7_15_g35182/U$3 ( \5143 , \5142 );
mnot \mul_7_15_g35182/U$4 ( \5144 , \4611 );
mor \mul_7_15_g35182/U$2 ( \5145 , \5143 , \5144 );
mnot \mul_7_15_fopt36302/U$1 ( \5146 , \4602 );
mnand \mul_7_15_g35307/U$1 ( \5147 , \4878 , \5146 );
mnand \mul_7_15_g35182/U$1 ( \5148 , \5145 , \5147 );
mnot \mul_7_15_g34795/U$4 ( \5149 , \5148 );
mor \mul_7_15_g34795/U$2 ( \5150 , \5136 , \5149 );
mor \mul_7_15_g34878/U$2 ( \5151 , \5148 , \5135 );
mnot \mul_7_15_g35681/U$3 ( \5152 , \4093 );
mnot \mul_7_15_g35681/U$4 ( \5153 , \4493 );
mor \mul_7_15_g35681/U$2 ( \5154 , \5152 , \5153 );
mnand \mul_7_15_g35853/U$1 ( \5155 , \4285 , \4349 );
mnand \mul_7_15_g35681/U$1 ( \5156 , \5154 , \5155 );
mnot \mul_7_15_g35185/U$3 ( \5157 , \5156 );
mnot \mul_7_15_g35185/U$4 ( \5158 , \4430 );
mor \mul_7_15_g35185/U$2 ( \5159 , \5157 , \5158 );
mbuf \mul_7_15_g35573/U$1 ( \5160 , \4800 );
mnand \mul_7_15_g35465/U$1 ( \5161 , \4891 , \5160 );
mnand \mul_7_15_g35185/U$1 ( \5162 , \5159 , \5161 );
mnand \mul_7_15_g34878/U$1 ( \5163 , \5151 , \5162 );
mnand \mul_7_15_g34795/U$1 ( \5164 , \5150 , \5163 );
mnot \mul_7_15_g34771/U$1 ( \5165 , \5164 );
mnot \mul_7_15_g34680/U$3 ( \5166 , \5165 );
mxor \mul_7_15_g36405/U$1 ( \5167 , \4870 , \4883 );
mxor \mul_7_15_g36405/U$1_r1 ( \5168 , \5167 , \4896 );
mnot \mul_7_15_g34680/U$4 ( \5169 , \5168 );
mor \mul_7_15_g34680/U$2 ( \5170 , \5166 , \5169 );
mnot \mul_7_15_g35635/U$3 ( \5171 , \4066 );
mnot \mul_7_15_g35635/U$4 ( \5172 , \4163 );
mor \mul_7_15_g35635/U$2 ( \5173 , \5171 , \5172 );
mnand \mul_7_15_g35803/U$1 ( \5174 , \4311 , \4519 );
mnand \mul_7_15_g35635/U$1 ( \5175 , \5173 , \5174 );
mnot \mul_7_15_g35193/U$3 ( \5176 , \5175 );
mnot \mul_7_15_g35193/U$4 ( \5177 , \4159 );
mor \mul_7_15_g35193/U$2 ( \5178 , \5176 , \5177 );
mnand \mul_7_15_g35327/U$1 ( \5179 , \4150 , \4908 );
mnand \mul_7_15_g35193/U$1 ( \5180 , \5178 , \5179 );
mnot \mul_7_15_g34786/U$3 ( \5181 , \5180 );
mnot \mul_7_15_g35714/U$3 ( \5182 , \4021 );
mnot \fopt36868/U$1 ( \5183 , \4110 );
mnot \mul_7_15_g35714/U$4 ( \5184 , \5183 );
mor \mul_7_15_g35714/U$2 ( \5185 , \5182 , \5184 );
mnand \mul_7_15_g35875/U$1 ( \5186 , \4106 , \4780 );
mnand \mul_7_15_g35714/U$1 ( \5187 , \5185 , \5186 );
mnot \mul_7_15_g35191/U$3 ( \5188 , \5187 );
mnot \mul_7_15_g35191/U$4 ( \5189 , \4710 );
mor \mul_7_15_g35191/U$2 ( \5190 , \5188 , \5189 );
mnand \mul_7_15_g35308/U$1 ( \5191 , \4957 , \4132 );
mnand \mul_7_15_g35191/U$1 ( \5192 , \5190 , \5191 );
mnot \mul_7_15_g34786/U$4 ( \5193 , \5192 );
mor \mul_7_15_g34786/U$2 ( \5194 , \5181 , \5193 );
mor \mul_7_15_g34873/U$2 ( \5195 , \5192 , \5180 );
mnot \mul_7_15_g35220/U$3 ( \5196 , \5122 );
mnot \mul_7_15_g35220/U$4 ( \5197 , \4632 );
mor \mul_7_15_g35220/U$2 ( \5198 , \5196 , \5197 );
mnand \mul_7_15_g36758/U$1 ( \5199 , \4453 , \4921 );
mnand \mul_7_15_g35220/U$1 ( \5200 , \5198 , \5199 );
mnand \mul_7_15_g34873/U$1 ( \5201 , \5195 , \5200 );
mnand \mul_7_15_g34786/U$1 ( \5202 , \5194 , \5201 );
mnand \mul_7_15_g34680/U$1 ( \5203 , \5170 , \5202 );
mnot \mul_7_15_g36385/U$2 ( \5204 , \5165 );
mnot \fopt36912/U$1 ( \5205 , \5168 );
mnand \mul_7_15_g36385/U$1 ( \5206 , \5204 , \5205 );
mand \mul_7_15_g36348/U$1 ( \5207 , \5203 , \5206 );
mxor \mul_7_15_g34449/U$1 ( \5208 , \5132 , \5207 );
mnot \mul_7_15_g34731/U$3 ( \5209 , \4982 );
mnot \mul_7_15_g34731/U$4 ( \5210 , \4978 );
mor \mul_7_15_g34731/U$2 ( \5211 , \5209 , \5210 );
mor \mul_7_15_g34731/U$5 ( \5212 , \4978 , \4982 );
mnand \mul_7_15_g34731/U$1 ( \5213 , \5211 , \5212 );
mnot \fopt36954/U$1 ( \5214 , \4996 );
mand \mul_7_15_g34648/U$2 ( \5215 , \5213 , \5214 );
mnot \mul_7_15_g34648/U$4 ( \5216 , \5213 );
mand \mul_7_15_g34648/U$3 ( \5217 , \5216 , \4996 );
mnor \mul_7_15_g34648/U$1 ( \5218 , \5215 , \5217 );
mxor \mul_7_15_g34449/U$1_r1 ( \5219 , \5208 , \5218 );
mxor \mul_7_15_g34322/U$1 ( \5220 , \5130 , \5219 );
mnot \mul_7_15_g35232/U$1 ( \5221 , \4951 );
mnot \mul_7_15_g34950/U$3 ( \5222 , \5221 );
mnot \mul_7_15_g34950/U$4 ( \5223 , \5100 );
mor \mul_7_15_g34950/U$2 ( \5224 , \5222 , \5223 );
mor \mul_7_15_g34950/U$5 ( \5225 , \5100 , \5221 );
mnand \mul_7_15_g34950/U$1 ( \5226 , \5224 , \5225 );
mnot \mul_7_15_g34918/U$1 ( \5227 , \5125 );
mand \mul_7_15_g34801/U$2 ( \5228 , \5226 , \5227 );
mnot \mul_7_15_g34801/U$4 ( \5229 , \5226 );
mand \mul_7_15_g34801/U$3 ( \5230 , \5229 , \5125 );
mnor \mul_7_15_g34801/U$1 ( \5231 , \5228 , \5230 );
mnot \mul_7_15_g34765/U$1 ( \5232 , \5231 );
mnot \g37169/U$3 ( \5233 , \5232 );
mbuf \fopt36914/U$1 ( \5234 , \5162 );
mand \mul_7_15_g34948/U$2 ( \5235 , \5148 , \5135 );
mnot \mul_7_15_g34948/U$4 ( \5236 , \5148 );
mand \mul_7_15_g34948/U$3 ( \5237 , \5236 , \5134 );
mnor \mul_7_15_g34948/U$1 ( \5238 , \5235 , \5237 );
mxor \mul_7_15_g36784/U$1 ( \5239 , \5234 , \5238 );
mnot \g37169/U$4 ( \5240 , \5239 );
mor \g37169/U$2 ( \5241 , \5233 , \5240 );
mnot \g37170/U$3 ( \5242 , \5231 );
mnot \mul_7_15_g34769/U$1 ( \5243 , \5239 );
mnot \g37170/U$4 ( \5244 , \5243 );
mor \g37170/U$2 ( \5245 , \5242 , \5244 );
mnor \mul_7_15_g34993/U$1 ( \5246 , \5124 , \5110 );
mnot \mul_7_15_g34939/U$2 ( \5247 , \5246 );
mnand \mul_7_15_g34939/U$1 ( \5248 , \5247 , \5125 );
mnot \mul_7_15_g35723/U$3 ( \5249 , \4026 );
mnot \mul_7_15_g35723/U$4 ( \5250 , \5183 );
mor \mul_7_15_g35723/U$2 ( \5251 , \5249 , \5250 );
mnand \mul_7_15_g35891/U$1 ( \5252 , \4106 , \4969 );
mnand \mul_7_15_g35723/U$1 ( \5253 , \5251 , \5252 );
mnot \mul_7_15_g35088/U$3 ( \5254 , \5253 );
mnot \mul_7_15_g35088/U$4 ( \5255 , \4129 );
mor \mul_7_15_g35088/U$2 ( \5256 , \5254 , \5255 );
mnand \mul_7_15_g35441/U$1 ( \5257 , \4133 , \5187 );
mnand \mul_7_15_g35088/U$1 ( \5258 , \5256 , \5257 );
mand \mul_7_15_g34868/U$1 ( \5259 , \5248 , \5258 );
mnand \g37170/U$1 ( \5260 , \5245 , \5259 );
mnand \g37169/U$1 ( \5261 , \5241 , \5260 );
mnot \mul_7_15_g34570/U$1 ( \5262 , \5261 );
mxor \mul_7_15_g34645/U$1 ( \5263 , \5164 , \5202 );
mxnor \mul_7_15_g34645/U$1_r1 ( \5264 , \5263 , \5205 );
mnand \mul_7_15_g34528/U$1 ( \5265 , \5262 , \5264 );
mbuf \mul_7_15_g35961/U$1 ( \5266 , \3241 );
mnot \mul_7_15_g36434/U$2 ( \5267 , \5266 );
mbuf \mul_7_15_fopt36327/U$1 ( \5268 , \3070 );
mnot \mul_7_15_g35898/U$2 ( \5269 , \5268 );
mnor \mul_7_15_g35898/U$1 ( \5270 , \5269 , \3241 );
mbuf \mul_7_15_g35897/U$1 ( \5271 , \5270 );
mnot \mul_7_15_g35896/U$1 ( \5272 , \5271 );
mnand \mul_7_15_g36434/U$1 ( \5273 , \5267 , \5272 );
mnot \mul_7_15_fopt36317/U$1 ( \5274 , \5268 );
mnot \mul_7_15_fopt36316/U$1 ( \5275 , \5274 );
mnand \mul_7_15_g35506/U$1 ( \5276 , \5273 , \5275 );
mnot \mul_7_15_g35265/U$2 ( \5277 , \5276 );
mnand \mul_7_15_g35770/U$1 ( \5278 , \4253 , \4079 );
mnand \mul_7_15_g35265/U$1 ( \5279 , \5277 , \5278 );
mnot \mul_7_15_g34953/U$3 ( \5280 , \5279 );
mnot \mul_7_15_g35609/U$3 ( \5281 , \4076 );
mnot \mul_7_15_g35609/U$4 ( \5282 , \4250 );
mor \mul_7_15_g35609/U$2 ( \5283 , \5281 , \5282 );
mnot \mul_7_15_g35946/U$1 ( \5284 , \4076 );
mnand \mul_7_15_g35879/U$1 ( \5285 , \5133 , \5284 );
mnand \mul_7_15_g35609/U$1 ( \5286 , \5283 , \5285 );
mnot \mul_7_15_g35059/U$3 ( \5287 , \5286 );
mnot \mul_7_15_g35059/U$4 ( \5288 , \4395 );
mor \mul_7_15_g35059/U$2 ( \5289 , \5287 , \5288 );
mnand \mul_7_15_g35252/U$1 ( \5290 , \5091 , \4200 );
mnand \mul_7_15_g35059/U$1 ( \5291 , \5289 , \5290 );
mnot \mul_7_15_g34953/U$4 ( \5292 , \5291 );
mor \mul_7_15_g34953/U$2 ( \5293 , \5280 , \5292 );
mnot \mul_7_15_g35514/U$1 ( \5294 , \5278 );
mnand \mul_7_15_g35264/U$1 ( \5295 , \5294 , \5276 );
mnand \mul_7_15_g34953/U$1 ( \5296 , \5293 , \5295 );
mnot \fopt36845/U$1 ( \5297 , \5296 );
mnot \mul_7_15_g34654/U$3 ( \5298 , \5297 );
mnot \mul_7_15_g35093/U$3 ( \5299 , \4611 );
mnot \mul_7_15_g35618/U$3 ( \5300 , \4094 );
mnot \mul_7_15_g36139/U$1 ( \5301 , \4616 );
mnot \mul_7_15_g35618/U$4 ( \5302 , \5301 );
mor \mul_7_15_g35618/U$2 ( \5303 , \5300 , \5302 );
mnand \mul_7_15_g37011/U$1 ( \5304 , \4616 , \4298 );
mnand \mul_7_15_g35618/U$1 ( \5305 , \5303 , \5304 );
mnot \mul_7_15_g35093/U$4 ( \5306 , \5305 );
mor \mul_7_15_g35093/U$2 ( \5307 , \5299 , \5306 );
mnand \mul_7_15_g35339/U$1 ( \5308 , \5142 , \4881 );
mnand \mul_7_15_g35093/U$1 ( \5309 , \5307 , \5308 );
mnot \mul_7_15_g34915/U$3 ( \5310 , \5309 );
mnot \mul_7_15_g35643/U$3 ( \5311 , \4017 );
mnot \mul_7_15_g35643/U$4 ( \5312 , \4163 );
mor \mul_7_15_g35643/U$2 ( \5313 , \5311 , \5312 );
mnand \mul_7_15_g35871/U$1 ( \5314 , \4164 , \4662 );
mnand \mul_7_15_g35643/U$1 ( \5315 , \5313 , \5314 );
mnot \mul_7_15_g35166/U$3 ( \5316 , \5315 );
mnot \mul_7_15_g35166/U$4 ( \5317 , \4159 );
mor \mul_7_15_g35166/U$2 ( \5318 , \5316 , \5317 );
mnand \mul_7_15_g35326/U$1 ( \5319 , \4317 , \5175 );
mnand \mul_7_15_g35166/U$1 ( \5320 , \5318 , \5319 );
mnot \mul_7_15_g34915/U$4 ( \5321 , \5320 );
mor \mul_7_15_g34915/U$2 ( \5322 , \5310 , \5321 );
mor \mul_7_15_g34937/U$2 ( \5323 , \5309 , \5320 );
mnot \mul_7_15_g35621/U$3 ( \5324 , \4095 );
mnot \mul_7_15_g35621/U$4 ( \5325 , \4332 );
mor \mul_7_15_g35621/U$2 ( \5326 , \5324 , \5325 );
mnand \mul_7_15_g35846/U$1 ( \5327 , \4283 , \4391 );
mnand \mul_7_15_g35621/U$1 ( \5328 , \5326 , \5327 );
mnot \mul_7_15_g35204/U$3 ( \5329 , \5328 );
mnot \mul_7_15_g35204/U$4 ( \5330 , \4430 );
mor \mul_7_15_g35204/U$2 ( \5331 , \5329 , \5330 );
mnand \mul_7_15_g35303/U$1 ( \5332 , \5156 , \4341 );
mnand \mul_7_15_g35204/U$1 ( \5333 , \5331 , \5332 );
mnand \mul_7_15_g34937/U$1 ( \5334 , \5323 , \5333 );
mnand \mul_7_15_g34915/U$1 ( \5335 , \5322 , \5334 );
mnot \mul_7_15_g34838/U$1 ( \5336 , \5335 );
mnot \mul_7_15_g34654/U$4 ( \5337 , \5336 );
mor \mul_7_15_g34654/U$2 ( \5338 , \5298 , \5337 );
mxor \g36942/U$1 ( \5339 , \5192 , \5180 );
mand \mul_7_15_g34859/U$2 ( \5340 , \5339 , \5200 );
mnot \mul_7_15_g34859/U$4 ( \5341 , \5339 );
mnot \fopt36934/U$1 ( \5342 , \5200 );
mand \mul_7_15_g34859/U$3 ( \5343 , \5341 , \5342 );
mnor \mul_7_15_g34859/U$1 ( \5344 , \5340 , \5343 );
mnand \mul_7_15_g34654/U$1 ( \5345 , \5338 , \5344 );
mnot \mul_7_15_g36393/U$2 ( \5346 , \5336 );
mbuf \fopt36844/U$1 ( \5347 , \5296 );
mnand \mul_7_15_g36393/U$1 ( \5348 , \5346 , \5347 );
mnand \mul_7_15_g34629/U$1 ( \5349 , \5345 , \5348 );
mbuf \fopt36936/U$1 ( \5350 , \5349 );
mand \mul_7_15_g34492/U$2 ( \5351 , \5265 , \5350 );
mnor \mul_7_15_g34527/U$1 ( \5352 , \5262 , \5264 );
mnor \mul_7_15_g34492/U$1 ( \5353 , \5351 , \5352 );
mxor \mul_7_15_g34322/U$1_r1 ( \5354 , \5220 , \5353 );
mxor \mul_7_15_g34501/U$1 ( \5355 , \5349 , \5264 );
mxnor \mul_7_15_g34501/U$1_r1 ( \5356 , \5355 , \5261 );
mnot \mul_7_15_g34475/U$1 ( \5357 , \5356 );
mnot \mul_7_15_g34694/U$3 ( \5358 , \5079 );
mnot \mul_7_15_g34766/U$1 ( \5359 , \5127 );
mnot \mul_7_15_g34694/U$4 ( \5360 , \5359 );
mor \mul_7_15_g34694/U$2 ( \5361 , \5358 , \5360 );
mnand \mul_7_15_g34713/U$1 ( \5362 , \5078 , \5127 );
mnand \mul_7_15_g34694/U$1 ( \5363 , \5361 , \5362 );
mnot \mul_7_15_g34756/U$1 ( \5364 , \5083 );
mand \mul_7_15_g34631/U$2 ( \5365 , \5363 , \5364 );
mnot \mul_7_15_g34631/U$4 ( \5366 , \5363 );
mand \mul_7_15_g34631/U$3 ( \5367 , \5366 , \5083 );
mnor \mul_7_15_g34631/U$1 ( \5368 , \5365 , \5367 );
mbuf \fopt37219/U$1 ( \5369 , \5368 );
mnot \fopt37218/U$1 ( \5370 , \5369 );
mnand \mul_7_15_g34435/U$1 ( \5371 , \5357 , \5370 );
mnot \mul_7_15_g35625/U$3 ( \5372 , \4198 );
mnot \mul_7_15_g35625/U$4 ( \5373 , \4935 );
mor \mul_7_15_g35625/U$2 ( \5374 , \5372 , \5373 );
mnand \mul_7_15_g35801/U$1 ( \5375 , \4934 , \4209 );
mnand \mul_7_15_g35625/U$1 ( \5376 , \5374 , \5375 );
mnot \mul_7_15_g35052/U$3 ( \5377 , \5376 );
mnot \mul_7_15_g35052/U$4 ( \5378 , \4944 );
mor \mul_7_15_g35052/U$2 ( \5379 , \5377 , \5378 );
mnand \mul_7_15_g35333/U$1 ( \5380 , \4863 , \5107 );
mnand \mul_7_15_g35052/U$1 ( \5381 , \5379 , \5380 );
mnot \mul_7_15_g34787/U$3 ( \5382 , \5381 );
mnot \mul_7_15_g35650/U$3 ( \5383 , \4072 );
mnot \mul_7_15_g35650/U$4 ( \5384 , \5183 );
mor \mul_7_15_g35650/U$2 ( \5385 , \5383 , \5384 );
mnand \mul_7_15_g35800/U$1 ( \5386 , \4110 , \5089 );
mnand \mul_7_15_g35650/U$1 ( \5387 , \5385 , \5386 );
mnot \mul_7_15_g35225/U$3 ( \5388 , \5387 );
mnot \mul_7_15_g35225/U$4 ( \5389 , \4128 );
mor \mul_7_15_g35225/U$2 ( \5390 , \5388 , \5389 );
mnand \mul_7_15_g35417/U$1 ( \5391 , \4132 , \5253 );
mnand \mul_7_15_g35225/U$1 ( \5392 , \5390 , \5391 );
mnot \mul_7_15_g35224/U$1 ( \5393 , \5392 );
mnot \mul_7_15_g35223/U$1 ( \5394 , \5393 );
mnot \mul_7_15_g34787/U$4 ( \5395 , \5394 );
mor \mul_7_15_g34787/U$2 ( \5396 , \5382 , \5395 );
mnot \mul_7_15_g35051/U$1 ( \5397 , \5381 );
mnot \mul_7_15_g34875/U$3 ( \5398 , \5397 );
mnot \mul_7_15_g34875/U$4 ( \5399 , \5393 );
mor \mul_7_15_g34875/U$2 ( \5400 , \5398 , \5399 );
mnot \mul_7_15_g35717/U$3 ( \5401 , \4780 );
mnot \mul_7_15_g35717/U$4 ( \5402 , \4311 );
mor \mul_7_15_g35717/U$2 ( \5403 , \5401 , \5402 );
mnand \mul_7_15_g35867/U$1 ( \5404 , \4163 , \4021 );
mnand \mul_7_15_g35717/U$1 ( \5405 , \5403 , \5404 );
mnot \mul_7_15_g35228/U$3 ( \5406 , \5405 );
mnot \mul_7_15_g35228/U$4 ( \5407 , \4159 );
mor \mul_7_15_g35228/U$2 ( \5408 , \5406 , \5407 );
mnand \mul_7_15_g35368/U$1 ( \5409 , \4317 , \5315 );
mnand \mul_7_15_g35228/U$1 ( \5410 , \5408 , \5409 );
mnand \mul_7_15_g34875/U$1 ( \5411 , \5400 , \5410 );
mnand \mul_7_15_g34787/U$1 ( \5412 , \5396 , \5411 );
mnot \mul_7_15_g34714/U$2 ( \5413 , \5412 );
mxor \mul_7_15_g34890/U$1 ( \5414 , \5276 , \5294 );
mxnor \mul_7_15_g34890/U$1_r1 ( \5415 , \5414 , \5291 );
mnand \mul_7_15_g34714/U$1 ( \5416 , \5413 , \5415 );
mnot \mul_7_15_g34563/U$3 ( \5417 , \5416 );
mnot \mul_7_15_g36021/U$1 ( \5418 , \4098 );
mnor \mul_7_15_g35899/U$1 ( \5419 , \4388 , \5418 );
mnot \mul_7_15_g35270/U$3 ( \5420 , \5271 );
mnot \mul_7_15_g35731/U$3 ( \5421 , \3997 );
mnot \mul_7_15_fopt36324/U$1 ( \5422 , \5268 );
mnot \mul_7_15_g35731/U$4 ( \5423 , \5422 );
mor \mul_7_15_g35731/U$2 ( \5424 , \5421 , \5423 );
mnot \mul_7_15_fopt36323/U$1 ( \5425 , \5422 );
mnand \mul_7_15_g35865/U$1 ( \5426 , \5425 , \4111 );
mnand \mul_7_15_g35731/U$1 ( \5427 , \5424 , \5426 );
mnot \mul_7_15_g35270/U$4 ( \5428 , \5427 );
mor \mul_7_15_g35270/U$2 ( \5429 , \5420 , \5428 );
mnot \mul_7_15_g35617/U$3 ( \5430 , \4051 );
mnot \mul_7_15_g35617/U$4 ( \5431 , \5422 );
mor \mul_7_15_g35617/U$2 ( \5432 , \5430 , \5431 );
mbuf \mul_7_15_fopt36313/U$1 ( \5433 , \5268 );
mnand \mul_7_15_g35787/U$1 ( \5434 , \5433 , \4135 );
mnand \mul_7_15_g35617/U$1 ( \5435 , \5432 , \5434 );
mnand \mul_7_15_g35306/U$1 ( \5436 , \5435 , \5266 );
mnand \mul_7_15_g35270/U$1 ( \5437 , \5429 , \5436 );
mxor \mul_7_15_g34815/U$4 ( \5438 , \5419 , \5437 );
mand \mul_7_15_g35667/U$2 ( \5439 , \4935 , \4094 );
mand \mul_7_15_g35667/U$3 ( \5440 , \4934 , \4298 );
mnor \mul_7_15_g35667/U$1 ( \5441 , \5439 , \5440 );
mor \mul_7_15_g35032/U$2 ( \5442 , \4943 , \5441 );
mnot \mul_7_15_g35624/U$1 ( \5443 , \5376 );
mor \mul_7_15_g35032/U$3 ( \5444 , \5443 , \4862 );
mnand \mul_7_15_g35032/U$1 ( \5445 , \5442 , \5444 );
mand \mul_7_15_g34815/U$3 ( \5446 , \5438 , \5445 );
mand \mul_7_15_g34815/U$5 ( \5447 , \5419 , \5437 );
mor \mul_7_15_g34815/U$2 ( \5448 , \5446 , \5447 );
mnot \mul_7_15_g35711/U$3 ( \5449 , \4969 );
mnot \mul_7_15_g35711/U$4 ( \5450 , \4311 );
mor \mul_7_15_g35711/U$2 ( \5451 , \5449 , \5450 );
mnand \mul_7_15_g36762/U$1 ( \5452 , \4163 , \4026 );
mnand \mul_7_15_g35711/U$1 ( \5453 , \5451 , \5452 );
mnot \mul_7_15_g35075/U$3 ( \5454 , \5453 );
mnot \mul_7_15_g35075/U$4 ( \5455 , \4158 );
mor \mul_7_15_g35075/U$2 ( \5456 , \5454 , \5455 );
mnand \mul_7_15_g35336/U$1 ( \5457 , \5405 , \4150 );
mnand \mul_7_15_g35075/U$1 ( \5458 , \5456 , \5457 );
mnot \mul_7_15_g34907/U$3 ( \5459 , \5458 );
mnot \mul_7_15_g35076/U$3 ( \5460 , \4610 );
mnot \mul_7_15_g35661/U$3 ( \5461 , \4097 );
mnot \mul_7_15_g35661/U$4 ( \5462 , \4746 );
mor \mul_7_15_g35661/U$2 ( \5463 , \5461 , \5462 );
mnand \mul_7_15_g35855/U$1 ( \5464 , \4745 , \4254 );
mnand \mul_7_15_g35661/U$1 ( \5465 , \5463 , \5464 );
mnot \mul_7_15_g35076/U$4 ( \5466 , \5465 );
mor \mul_7_15_g35076/U$2 ( \5467 , \5460 , \5466 );
mnot \mul_7_15_g35724/U$3 ( \5468 , \4096 );
mnot \mul_7_15_g35724/U$4 ( \5469 , \5138 );
mor \mul_7_15_g35724/U$2 ( \5470 , \5468 , \5469 );
mnand \mul_7_15_g35828/U$1 ( \5471 , \4615 , \4372 );
mnand \mul_7_15_g35724/U$1 ( \5472 , \5470 , \5471 );
mnand \mul_7_15_g35359/U$1 ( \5473 , \4754 , \5472 );
mnand \mul_7_15_g35076/U$1 ( \5474 , \5467 , \5473 );
mnot \mul_7_15_g34907/U$4 ( \5475 , \5474 );
mor \mul_7_15_g34907/U$2 ( \5476 , \5459 , \5475 );
mor \mul_7_15_g34931/U$2 ( \5477 , \5474 , \5458 );
mnot \mul_7_15_g35692/U$3 ( \5478 , \4076 );
mnot \mul_7_15_g35692/U$4 ( \5479 , \4134 );
mor \mul_7_15_g35692/U$2 ( \5480 , \5478 , \5479 );
mnand \mul_7_15_g35863/U$1 ( \5481 , \4106 , \5284 );
mnand \mul_7_15_g35692/U$1 ( \5482 , \5480 , \5481 );
mnot \mul_7_15_g35197/U$3 ( \5483 , \5482 );
mnot \mul_7_15_g35197/U$4 ( \5484 , \4710 );
mor \mul_7_15_g35197/U$2 ( \5485 , \5483 , \5484 );
mnand \mul_7_15_g35370/U$1 ( \5486 , \5387 , \4132 );
mnand \mul_7_15_g35197/U$1 ( \5487 , \5485 , \5486 );
mnand \mul_7_15_g34931/U$1 ( \5488 , \5477 , \5487 );
mnand \mul_7_15_g34907/U$1 ( \5489 , \5476 , \5488 );
mxor \mul_7_15_g34637/U$4 ( \5490 , \5448 , \5489 );
mnot \mul_7_15_g35701/U$3 ( \5491 , \4017 );
mnot \mul_7_15_g35701/U$4 ( \5492 , \4332 );
mor \mul_7_15_g35701/U$2 ( \5493 , \5491 , \5492 );
mnand \mul_7_15_g35833/U$1 ( \5494 , \4283 , \4662 );
mnand \mul_7_15_g35701/U$1 ( \5495 , \5493 , \5494 );
mnot \mul_7_15_g35181/U$3 ( \5496 , \5495 );
mnot \fopt/U$1 ( \5497 , \4278 );
mnot \mul_7_15_g35181/U$4 ( \5498 , \5497 );
mor \mul_7_15_g35181/U$2 ( \5499 , \5496 , \5498 );
mnot \mul_7_15_g35718/U$3 ( \5500 , \4066 );
mnot \mul_7_15_g35718/U$4 ( \5501 , \4493 );
mor \mul_7_15_g35718/U$2 ( \5502 , \5500 , \5501 );
mnand \mul_7_15_g35848/U$1 ( \5503 , \4283 , \4519 );
mnand \mul_7_15_g35718/U$1 ( \5504 , \5502 , \5503 );
mnand \mul_7_15_g35330/U$1 ( \5505 , \5504 , \4800 );
mnand \mul_7_15_g35181/U$1 ( \5506 , \5499 , \5505 );
mnot \mul_7_15_g35074/U$3 ( \5507 , \4449 );
mnot \mul_7_15_g35644/U$3 ( \5508 , \4095 );
mnot \mul_7_15_g35644/U$4 ( \5509 , \5112 );
mor \mul_7_15_g35644/U$2 ( \5510 , \5508 , \5509 );
mnand \mul_7_15_g35827/U$1 ( \5511 , \4536 , \4391 );
mnand \mul_7_15_g35644/U$1 ( \5512 , \5510 , \5511 );
mnot \mul_7_15_g35074/U$4 ( \5513 , \5512 );
mor \mul_7_15_g35074/U$2 ( \5514 , \5507 , \5513 );
mnot \mul_7_15_g35636/U$3 ( \5515 , \4093 );
mnot \mul_7_15_g35636/U$4 ( \5516 , \5112 );
mor \mul_7_15_g35636/U$2 ( \5517 , \5515 , \5516 );
mnand \mul_7_15_g35851/U$1 ( \5518 , \4729 , \4349 );
mnand \mul_7_15_g35636/U$1 ( \5519 , \5517 , \5518 );
mnand \mul_7_15_g35332/U$1 ( \5520 , \5519 , \4452 );
mnand \mul_7_15_g35074/U$1 ( \5521 , \5514 , \5520 );
mxor \mul_7_15_g34804/U$4 ( \5522 , \5506 , \5521 );
mnot \mul_7_15_g35599/U$3 ( \5523 , \4082 );
mnot \mul_7_15_g35599/U$4 ( \5524 , \4388 );
mor \mul_7_15_g35599/U$2 ( \5525 , \5523 , \5524 );
mnot \mul_7_15_g36150/U$1 ( \5526 , \4082 );
mnand \mul_7_15_g35844/U$1 ( \5527 , \4100 , \5526 );
mnand \mul_7_15_g35599/U$1 ( \5528 , \5525 , \5527 );
mnot \mul_7_15_g35053/U$3 ( \5529 , \5528 );
mnot \mul_7_15_g35053/U$4 ( \5530 , \4395 );
mor \mul_7_15_g35053/U$2 ( \5531 , \5529 , \5530 );
mnot \mul_7_15_g35605/U$3 ( \5532 , \4079 );
mnot \mul_7_15_g35605/U$4 ( \5533 , \4101 );
mor \mul_7_15_g35605/U$2 ( \5534 , \5532 , \5533 );
mnot \mul_7_15_g36131/U$1 ( \5535 , \4079 );
mnand \mul_7_15_g35868/U$1 ( \5536 , \4100 , \5535 );
mnand \mul_7_15_g35605/U$1 ( \5537 , \5534 , \5536 );
mnand \mul_7_15_g35250/U$1 ( \5538 , \5537 , \4200 );
mnand \mul_7_15_g35053/U$1 ( \5539 , \5531 , \5538 );
mand \mul_7_15_g34804/U$3 ( \5540 , \5522 , \5539 );
mand \mul_7_15_g34804/U$5 ( \5541 , \5506 , \5521 );
mor \mul_7_15_g34804/U$2 ( \5542 , \5540 , \5541 );
mand \mul_7_15_g34637/U$3 ( \5543 , \5490 , \5542 );
mand \mul_7_15_g34637/U$5 ( \5544 , \5448 , \5489 );
mor \mul_7_15_g34637/U$2 ( \5545 , \5543 , \5544 );
mnot \mul_7_15_g34563/U$4 ( \5546 , \5545 );
mor \mul_7_15_g34563/U$2 ( \5547 , \5417 , \5546 );
mnot \mul_7_15_g36392/U$2 ( \5548 , \5415 );
mnand \mul_7_15_g36392/U$1 ( \5549 , \5548 , \5412 );
mnand \mul_7_15_g34563/U$1 ( \5550 , \5547 , \5549 );
mnot \mul_7_15_g34472/U$3 ( \5551 , \5550 );
mand \g37272/U$2 ( \5552 , \5296 , \5336 );
mnot \g37272/U$4 ( \5553 , \5296 );
mand \g37272/U$3 ( \5554 , \5553 , \5335 );
mor \g37272/U$1 ( \5555 , \5552 , \5554 );
mand \mul_7_15_g34649/U$2 ( \5556 , \5555 , \5344 );
mnot \mul_7_15_g34649/U$4 ( \5557 , \5555 );
mnot \mul_7_15_g34758/U$1 ( \5558 , \5344 );
mand \mul_7_15_g34649/U$3 ( \5559 , \5557 , \5558 );
mnor \mul_7_15_g34649/U$1 ( \5560 , \5556 , \5559 );
mnot \mul_7_15_fopt36213/U$1 ( \5561 , \5560 );
mnot \mul_7_15_g35302/U$3 ( \5562 , \5435 );
mnot \mul_7_15_g35302/U$4 ( \5563 , \5271 );
mor \mul_7_15_g35302/U$2 ( \5564 , \5562 , \5563 );
mnand \mul_7_15_g35786/U$1 ( \5565 , \5275 , \5266 );
mnand \mul_7_15_g35302/U$1 ( \5566 , \5564 , \5565 );
mnot \mul_7_15_g35216/U$3 ( \5567 , \5504 );
mnot \mul_7_15_g35216/U$4 ( \5568 , \4797 );
mor \mul_7_15_g35216/U$2 ( \5569 , \5567 , \5568 );
mnand \mul_7_15_g36427/U$1 ( \5570 , \5328 , \4800 );
mnand \mul_7_15_g35216/U$1 ( \5571 , \5569 , \5570 );
mxor \mul_7_15_g34836/U$4 ( \5572 , \5566 , \5571 );
mnot \mul_7_15_g35215/U$3 ( \5573 , \5472 );
mnot \mul_7_15_g35215/U$4 ( \5574 , \4611 );
mor \mul_7_15_g35215/U$2 ( \5575 , \5573 , \5574 );
mnand \mul_7_15_g35363/U$1 ( \5576 , \5305 , \4881 );
mnand \mul_7_15_g35215/U$1 ( \5577 , \5575 , \5576 );
mand \mul_7_15_g34836/U$3 ( \5578 , \5572 , \5577 );
mand \mul_7_15_g34836/U$5 ( \5579 , \5566 , \5571 );
mor \mul_7_15_g34836/U$2 ( \5580 , \5578 , \5579 );
mnot \mul_7_15_g34691/U$3 ( \5581 , \5580 );
mxor \mul_7_15_g36767/U$1 ( \5582 , \5309 , \5320 );
mxor \mul_7_15_g36767/U$1_r1 ( \5583 , \5582 , \5333 );
mnot \mul_7_15_g34691/U$4 ( \5584 , \5583 );
mor \mul_7_15_g34691/U$2 ( \5585 , \5581 , \5584 );
mor \mul_7_15_g34721/U$2 ( \5586 , \5583 , \5580 );
mand \mul_7_15_g35771/U$1 ( \5587 , \4100 , \4082 );
mnot \mul_7_15_g34929/U$3 ( \5588 , \5587 );
mnot \mul_7_15_g35071/U$3 ( \5589 , \5537 );
mnot \mul_7_15_g35071/U$4 ( \5590 , \4395 );
mor \mul_7_15_g35071/U$2 ( \5591 , \5589 , \5590 );
mnand \mul_7_15_g35262/U$1 ( \5592 , \5286 , \4200 );
mnand \mul_7_15_g35071/U$1 ( \5593 , \5591 , \5592 );
mnot \mul_7_15_g34929/U$4 ( \5594 , \5593 );
mor \mul_7_15_g34929/U$2 ( \5595 , \5588 , \5594 );
mor \mul_7_15_g34942/U$2 ( \5596 , \5593 , \5587 );
mnot \mul_7_15_g35222/U$3 ( \5597 , \4449 );
mnot \mul_7_15_g35222/U$4 ( \5598 , \5519 );
mor \mul_7_15_g35222/U$2 ( \5599 , \5597 , \5598 );
mnand \mul_7_15_g35429/U$1 ( \5600 , \4452 , \5116 );
mnand \mul_7_15_g35222/U$1 ( \5601 , \5599 , \5600 );
mnand \mul_7_15_g34942/U$1 ( \5602 , \5596 , \5601 );
mnand \mul_7_15_g34929/U$1 ( \5603 , \5595 , \5602 );
mnand \mul_7_15_g34721/U$1 ( \5604 , \5586 , \5603 );
mnand \mul_7_15_g34691/U$1 ( \5605 , \5585 , \5604 );
mnot \mul_7_15_g34635/U$1 ( \5606 , \5605 );
mnand \mul_7_15_g34552/U$1 ( \5607 , \5561 , \5606 );
mnot \mul_7_15_g34472/U$4 ( \5608 , \5607 );
mor \mul_7_15_g34472/U$2 ( \5609 , \5551 , \5608 );
mnot \mul_7_15_g36334/U$2 ( \5610 , \5561 );
mnand \mul_7_15_g36334/U$1 ( \5611 , \5610 , \5605 );
mnand \mul_7_15_g34472/U$1 ( \5612 , \5609 , \5611 );
mbuf \mul_7_15_g34450/U$1 ( \5613 , \5612 );
mand \mul_7_15_g34368/U$2 ( \5614 , \5371 , \5613 );
mnot \fopt37217/U$1 ( \5615 , \5369 );
mnor \mul_7_15_g34446/U$1 ( \5616 , \5357 , \5615 );
mnor \mul_7_15_g34368/U$1 ( \5617 , \5614 , \5616 );
mnand \mul_7_15_g34284/U$1 ( \5618 , \5354 , \5617 );
mxor \mul_7_15_g34322/U$4 ( \5619 , \5130 , \5219 );
mand \mul_7_15_g34322/U$3 ( \5620 , \5619 , \5353 );
mand \mul_7_15_g34322/U$5 ( \5621 , \5130 , \5219 );
mor \mul_7_15_g34322/U$2 ( \5622 , \5620 , \5621 );
mnot \mul_7_15_g34730/U$3 ( \5623 , \4807 );
mnot \mul_7_15_g34730/U$4 ( \5624 , \4773 );
mor \mul_7_15_g34730/U$2 ( \5625 , \5623 , \5624 );
mnand \mul_7_15_g34740/U$1 ( \5626 , \4804 , \4772 );
mnand \mul_7_15_g34730/U$1 ( \5627 , \5625 , \5626 );
mnot \mul_7_15_g34839/U$1 ( \5628 , \4812 );
mand \mul_7_15_g34647/U$2 ( \5629 , \5627 , \5628 );
mnot \mul_7_15_g34647/U$4 ( \5630 , \5627 );
mand \mul_7_15_g34647/U$3 ( \5631 , \5630 , \4812 );
mnor \mul_7_15_g34647/U$1 ( \5632 , \5629 , \5631 );
mxor \mul_7_15_g34457/U$1 ( \5633 , \4847 , \4930 );
mxnor \mul_7_15_g34457/U$1_r1 ( \5634 , \5633 , \4999 );
mxor \mul_7_15_g34298/U$1 ( \5635 , \5632 , \5634 );
mxor \mul_7_15_g34449/U$4 ( \5636 , \5132 , \5207 );
mand \mul_7_15_g34449/U$3 ( \5637 , \5636 , \5218 );
mand \mul_7_15_g34449/U$5 ( \5638 , \5132 , \5207 );
mor \mul_7_15_g34449/U$2 ( \5639 , \5637 , \5638 );
mxor \mul_7_15_g34298/U$1_r1 ( \5640 , \5635 , \5639 );
mnand \mul_7_15_g34274/U$1 ( \5641 , \5622 , \5640 );
mxor \mul_7_15_g34298/U$4 ( \5642 , \5632 , \5634 );
mand \mul_7_15_g34298/U$3 ( \5643 , \5642 , \5639 );
mand \mul_7_15_g34298/U$5 ( \5644 , \5632 , \5634 );
mor \mul_7_15_g34298/U$2 ( \5645 , \5643 , \5644 );
mxor \mul_7_15_g34394/U$1 ( \5646 , \4837 , \5001 );
mxnor \mul_7_15_g34394/U$1_r1 ( \5647 , \5646 , \4834 );
mnand \mul_7_15_g34271/U$1 ( \5648 , \5645 , \5647 );
mand \mul_7_15_g34235/U$1 ( \5649 , \5618 , \5641 , \5648 );
mxor \mul_7_15_g34376/U$1 ( \5650 , \5368 , \5612 );
mxnor \mul_7_15_g34376/U$1_r1 ( \5651 , \5650 , \5356 );
mxor \mul_7_15_g34581/U$1 ( \5652 , \5239 , \5232 );
mxnor \mul_7_15_g34581/U$1_r1 ( \5653 , \5652 , \5259 );
mxor \mul_7_15_g34675/U$1 ( \5654 , \5580 , \5603 );
mxnor \mul_7_15_g34675/U$1_r1 ( \5655 , \5654 , \5583 );
mnot \mul_7_15_g34788/U$3 ( \5656 , \5248 );
mnot \mul_7_15_g35087/U$1 ( \5657 , \5258 );
mnot \mul_7_15_g34788/U$4 ( \5658 , \5657 );
mand \mul_7_15_g34788/U$2 ( \5659 , \5656 , \5658 );
mand \mul_7_15_g34788/U$5 ( \5660 , \5248 , \5657 );
mnor \mul_7_15_g34788/U$1 ( \5661 , \5659 , \5660 );
mbuf \mul_7_15_g34768/U$1 ( \5662 , \5661 );
mnand \mul_7_15_g34573/U$1 ( \5663 , \5655 , \5662 );
mxor \mul_7_15_g34836/U$1 ( \5664 , \5566 , \5571 );
mxor \mul_7_15_g34836/U$1_r1 ( \5665 , \5664 , \5577 );
mnot \mul_7_15_g34689/U$3 ( \5666 , \5665 );
mxor \mul_7_15_g34901/U$1 ( \5667 , \5587 , \5601 );
mxnor \mul_7_15_g34901/U$1_r1 ( \5668 , \5667 , \5593 );
mnot \mul_7_15_g34824/U$1 ( \5669 , \5668 );
mnot \mul_7_15_g34689/U$4 ( \5670 , \5669 );
mor \mul_7_15_g34689/U$2 ( \5671 , \5666 , \5670 );
mnot \mul_7_15_g34716/U$3 ( \5672 , \5668 );
mnot \mul_7_15_g34834/U$1 ( \5673 , \5665 );
mnot \mul_7_15_g34716/U$4 ( \5674 , \5673 );
mor \mul_7_15_g34716/U$2 ( \5675 , \5672 , \5674 );
mnot \mul_7_15_g34967/U$3 ( \5676 , \5397 );
mnot \mul_7_15_g34967/U$4 ( \5677 , \5392 );
mor \mul_7_15_g34967/U$2 ( \5678 , \5676 , \5677 );
mor \mul_7_15_g34967/U$5 ( \5679 , \5397 , \5392 );
mnand \mul_7_15_g34967/U$1 ( \5680 , \5678 , \5679 );
mnot \mul_7_15_g35227/U$1 ( \5681 , \5410 );
mand \mul_7_15_g34857/U$2 ( \5682 , \5680 , \5681 );
mnot \mul_7_15_g34857/U$4 ( \5683 , \5680 );
mand \mul_7_15_g34857/U$3 ( \5684 , \5683 , \5410 );
mnor \mul_7_15_g34857/U$1 ( \5685 , \5682 , \5684 );
mnot \fopt36856/U$1 ( \5686 , \5685 );
mnand \mul_7_15_g34716/U$1 ( \5687 , \5675 , \5686 );
mnand \mul_7_15_g34689/U$1 ( \5688 , \5671 , \5687 );
mand \mul_7_15_g34531/U$2 ( \5689 , \5663 , \5688 );
mnor \mul_7_15_g34572/U$1 ( \5690 , \5655 , \5662 );
mnor \mul_7_15_g34531/U$1 ( \5691 , \5689 , \5690 );
mxor \mul_7_15_g34373/U$4 ( \5692 , \5653 , \5691 );
mnot \mul_7_15_g34549/U$3 ( \5693 , \5605 );
mnot \mul_7_15_g34549/U$4 ( \5694 , \5561 );
mor \mul_7_15_g34549/U$2 ( \5695 , \5693 , \5694 );
mnand \mul_7_15_g34553/U$1 ( \5696 , \5606 , \5560 );
mnand \mul_7_15_g34549/U$1 ( \5697 , \5695 , \5696 );
mnot \mul_7_15_g34544/U$1 ( \5698 , \5550 );
mand \mul_7_15_g34482/U$2 ( \5699 , \5697 , \5698 );
mnot \mul_7_15_g34482/U$4 ( \5700 , \5697 );
mand \mul_7_15_g34482/U$3 ( \5701 , \5700 , \5550 );
mnor \mul_7_15_g34482/U$1 ( \5702 , \5699 , \5701 );
mand \mul_7_15_g34373/U$3 ( \5703 , \5692 , \5702 );
mand \mul_7_15_g34373/U$5 ( \5704 , \5653 , \5691 );
mor \mul_7_15_g34373/U$2 ( \5705 , \5703 , \5704 );
mnand \mul_7_15_g34306/U$1 ( \5706 , \5651 , \5705 );
mand \mul_7_15_g34216/U$1 ( \5707 , \5649 , \5706 );
mnot \mul_7_15_g34493/U$3 ( \5708 , \5655 );
mnot \mul_7_15_g34535/U$3 ( \5709 , \5661 );
mnot \mul_7_15_g34535/U$4 ( \5710 , \5688 );
mor \mul_7_15_g34535/U$2 ( \5711 , \5709 , \5710 );
mor \mul_7_15_g34535/U$5 ( \5712 , \5661 , \5688 );
mnand \mul_7_15_g34535/U$1 ( \5713 , \5711 , \5712 );
mnot \mul_7_15_g34493/U$4 ( \5714 , \5713 );
mor \mul_7_15_g34493/U$2 ( \5715 , \5708 , \5714 );
mor \mul_7_15_g34493/U$5 ( \5716 , \5655 , \5713 );
mnand \mul_7_15_g34493/U$1 ( \5717 , \5715 , \5716 );
mnot \mul_7_15_g34476/U$1 ( \5718 , \5717 );
mnot \mul_7_15_g34393/U$3 ( \5719 , \5718 );
mxor \g37229/U$1 ( \5720 , \5412 , \5415 );
mxnor \g37229/U$1_r1 ( \5721 , \5720 , \5545 );
mnot \mul_7_15_g34434/U$3 ( \5722 , \5721 );
mxor \mul_7_15_g34637/U$1 ( \5723 , \5448 , \5489 );
mxor \mul_7_15_g34637/U$1_r1 ( \5724 , \5723 , \5542 );
mnot \mul_7_15_g34636/U$1 ( \5725 , \5724 );
mnot \mul_7_15_g35522/U$3 ( \5726 , \5418 );
mnot \mul_7_15_g35522/U$4 ( \5727 , \4182 );
mor \mul_7_15_g35522/U$2 ( \5728 , \5726 , \5727 );
mnand \mul_7_15_g35522/U$1 ( \5729 , \5728 , \4110 );
mnot \mul_7_15_g36432/U$2 ( \5730 , \4182 );
mnand \mul_7_15_g36432/U$1 ( \5731 , \5730 , \4098 );
mnand \mul_7_15_g35493/U$1 ( \5732 , \4102 , \5729 , \5731 );
mnot \mul_7_15_g35715/U$3 ( \5733 , \4096 );
mnot \mul_7_15_g35715/U$4 ( \5734 , \4935 );
mor \mul_7_15_g35715/U$2 ( \5735 , \5733 , \5734 );
mnand \mul_7_15_g35876/U$1 ( \5736 , \2945 , \4372 );
mnand \mul_7_15_g35715/U$1 ( \5737 , \5735 , \5736 );
mnot \mul_7_15_g35043/U$3 ( \5738 , \5737 );
mnot \mul_7_15_g35043/U$4 ( \5739 , \4944 );
mor \mul_7_15_g35043/U$2 ( \5740 , \5738 , \5739 );
mnot \mul_7_15_g35331/U$2 ( \5741 , \5441 );
mnand \mul_7_15_g35331/U$1 ( \5742 , \5741 , \4863 );
mnand \mul_7_15_g35043/U$1 ( \5743 , \5740 , \5742 );
mnot \mul_7_15_g35042/U$1 ( \5744 , \5743 );
mnor \mul_7_15_g35004/U$1 ( \5745 , \5732 , \5744 );
mxor \mul_7_15_g34815/U$1 ( \5746 , \5419 , \5437 );
mxor \mul_7_15_g34815/U$1_r1 ( \5747 , \5746 , \5445 );
mxor \mul_7_15_g34643/U$4 ( \5748 , \5745 , \5747 );
mnot \mul_7_15_g35743/U$3 ( \5749 , \4198 );
mnot \mul_7_15_g35743/U$4 ( \5750 , \5422 );
mor \mul_7_15_g35743/U$2 ( \5751 , \5749 , \5750 );
mnand \mul_7_15_g35815/U$1 ( \5752 , \5433 , \4209 );
mnand \mul_7_15_g35743/U$1 ( \5753 , \5751 , \5752 );
mnot \mul_7_15_g35289/U$3 ( \5754 , \5753 );
mnot \mul_7_15_g35289/U$4 ( \5755 , \5271 );
mor \mul_7_15_g35289/U$2 ( \5756 , \5754 , \5755 );
mnand \mul_7_15_g35343/U$1 ( \5757 , \5427 , \5266 );
mnand \mul_7_15_g35289/U$1 ( \5758 , \5756 , \5757 );
mnot \mul_7_15_g35744/U$3 ( \5759 , \4098 );
mnot \mul_7_15_g35744/U$4 ( \5760 , \4346 );
mor \mul_7_15_g35744/U$2 ( \5761 , \5759 , \5760 );
mnand \mul_7_15_g35902/U$1 ( \5762 , \4100 , \5418 );
mnand \mul_7_15_g35744/U$1 ( \5763 , \5761 , \5762 );
mnot \mul_7_15_g35067/U$3 ( \5764 , \5763 );
mnot \mul_7_15_g35067/U$4 ( \5765 , \4194 );
mor \mul_7_15_g35067/U$2 ( \5766 , \5764 , \5765 );
mnand \mul_7_15_g35257/U$1 ( \5767 , \5528 , \4200 );
mnand \mul_7_15_g35067/U$1 ( \5768 , \5766 , \5767 );
mxor \mul_7_15_g34767/U$4 ( \5769 , \5758 , \5768 );
mand \mul_7_15_g35694/U$2 ( \5770 , \4519 , \4458 );
mnot \mul_7_15_g35694/U$4 ( \5771 , \4519 );
mand \mul_7_15_g35694/U$3 ( \5772 , \5771 , \4535 );
mnor \mul_7_15_g35694/U$1 ( \5773 , \5770 , \5772 );
mnot \mul_7_15_g35693/U$1 ( \5774 , \5773 );
mnot \mul_7_15_g35133/U$3 ( \5775 , \5774 );
mnot \mul_7_15_g35133/U$4 ( \5776 , \4632 );
mor \mul_7_15_g35133/U$2 ( \5777 , \5775 , \5776 );
mnand \mul_7_15_g35350/U$1 ( \5778 , \4453 , \5512 );
mnand \mul_7_15_g35133/U$1 ( \5779 , \5777 , \5778 );
mand \mul_7_15_g34767/U$3 ( \5780 , \5769 , \5779 );
mand \mul_7_15_g34767/U$5 ( \5781 , \5758 , \5768 );
mor \mul_7_15_g34767/U$2 ( \5782 , \5780 , \5781 );
mand \mul_7_15_g34643/U$3 ( \5783 , \5748 , \5782 );
mand \mul_7_15_g34643/U$5 ( \5784 , \5745 , \5747 );
mor \mul_7_15_g34643/U$2 ( \5785 , \5783 , \5784 );
mnot \mul_7_15_g34642/U$1 ( \5786 , \5785 );
mnand \mul_7_15_g34576/U$1 ( \5787 , \5725 , \5786 );
mxor \mul_7_15_g34804/U$1 ( \5788 , \5506 , \5521 );
mxor \mul_7_15_g34804/U$1_r1 ( \5789 , \5788 , \5539 );
mnot \mul_7_15_g34690/U$3 ( \5790 , \5789 );
mnot \mul_7_15_g35721/U$3 ( \5791 , \4093 );
mnot \mul_7_15_g35721/U$4 ( \5792 , \4746 );
mor \mul_7_15_g35721/U$2 ( \5793 , \5791 , \5792 );
mnand \mul_7_15_g35798/U$1 ( \5794 , \4615 , \4349 );
mnand \mul_7_15_g35721/U$1 ( \5795 , \5793 , \5794 );
mnot \mul_7_15_g35200/U$3 ( \5796 , \5795 );
mnot \mul_7_15_g35200/U$4 ( \5797 , \4610 );
mor \mul_7_15_g35200/U$2 ( \5798 , \5796 , \5797 );
mnand \mul_7_15_g35425/U$1 ( \5799 , \5465 , \5146 );
mnand \mul_7_15_g35200/U$1 ( \5800 , \5798 , \5799 );
mbuf \fopt36703/U$1 ( \5801 , \5800 );
mnot \mul_7_15_g34908/U$3 ( \5802 , \5801 );
mnot \fopt36886/U$1 ( \5803 , \4158 );
mnot \mul_7_15_g35175/U$3 ( \5804 , \5803 );
mand \mul_7_15_g35709/U$2 ( \5805 , \5089 , \4170 );
mnot \mul_7_15_g35709/U$4 ( \5806 , \5089 );
mand \mul_7_15_g35709/U$3 ( \5807 , \5806 , \4163 );
mnor \mul_7_15_g35709/U$1 ( \5808 , \5805 , \5807 );
mnot \mul_7_15_g35175/U$4 ( \5809 , \5808 );
mand \mul_7_15_g35175/U$2 ( \5810 , \5804 , \5809 );
mnot \mul_7_15_g36430/U$2 ( \5811 , \5453 );
mnor \mul_7_15_g36430/U$1 ( \5812 , \5811 , \4151 );
mnor \mul_7_15_g35175/U$1 ( \5813 , \5810 , \5812 );
mnot \mul_7_15_g35174/U$1 ( \5814 , \5813 );
mnot \mul_7_15_g34908/U$4 ( \5815 , \5814 );
mor \mul_7_15_g34908/U$2 ( \5816 , \5802 , \5815 );
mor \mul_7_15_g34932/U$2 ( \5817 , \5814 , \5801 );
mnot \g37140/U$3 ( \5818 , \4278 );
mand \mul_7_15_g35690/U$2 ( \5819 , \4021 , \4332 );
mnot \mul_7_15_g35690/U$4 ( \5820 , \4021 );
mand \mul_7_15_g35690/U$3 ( \5821 , \5820 , \4283 );
mnor \mul_7_15_g35690/U$1 ( \5822 , \5819 , \5821 );
mnot \g37140/U$4 ( \5823 , \5822 );
mand \g37140/U$2 ( \5824 , \5818 , \5823 );
mand \g37140/U$5 ( \5825 , \5495 , \4266 );
mnor \g37140/U$1 ( \5826 , \5824 , \5825 );
mnot \fopt36712/U$1 ( \5827 , \5826 );
mnand \mul_7_15_g34932/U$1 ( \5828 , \5817 , \5827 );
mnand \mul_7_15_g34908/U$1 ( \5829 , \5816 , \5828 );
mnot \mul_7_15_g34690/U$4 ( \5830 , \5829 );
mor \mul_7_15_g34690/U$2 ( \5831 , \5790 , \5830 );
mor \mul_7_15_g34717/U$2 ( \5832 , \5789 , \5829 );
mxor \mul_7_15_g36413/U$1 ( \5833 , \5474 , \5458 );
mxnor \mul_7_15_g36413/U$1_r1 ( \5834 , \5833 , \5487 );
mnot \mul_7_15_g34840/U$1 ( \5835 , \5834 );
mnand \mul_7_15_g34717/U$1 ( \5836 , \5832 , \5835 );
mnand \mul_7_15_g34690/U$1 ( \5837 , \5831 , \5836 );
mand \mul_7_15_g34490/U$2 ( \5838 , \5787 , \5837 );
mand \mul_7_15_g34545/U$2 ( \5839 , \5785 , \5724 );
mnor \mul_7_15_g34490/U$1 ( \5840 , \5838 , \5839 );
mnot \mul_7_15_g34434/U$4 ( \5841 , \5840 );
mor \mul_7_15_g34434/U$2 ( \5842 , \5722 , \5841 );
mor \mul_7_15_g34434/U$5 ( \5843 , \5721 , \5840 );
mnand \mul_7_15_g34434/U$1 ( \5844 , \5842 , \5843 );
mnot \mul_7_15_g34393/U$4 ( \5845 , \5844 );
mor \mul_7_15_g34393/U$2 ( \5846 , \5719 , \5845 );
mnot \mul_7_15_g34477/U$1 ( \5847 , \5717 );
mor \mul_7_15_g34393/U$5 ( \5848 , \5847 , \5844 );
mnand \mul_7_15_g34393/U$1 ( \5849 , \5846 , \5848 );
mnot \mul_7_15_g34700/U$3 ( \5850 , \5665 );
mnot \mul_7_15_g34700/U$4 ( \5851 , \5685 );
mor \mul_7_15_g34700/U$2 ( \5852 , \5850 , \5851 );
mor \mul_7_15_g34700/U$5 ( \5853 , \5665 , \5685 );
mnand \mul_7_15_g34700/U$1 ( \5854 , \5852 , \5853 );
mand \mul_7_15_g34644/U$2 ( \5855 , \5854 , \5669 );
mnot \mul_7_15_g34644/U$4 ( \5856 , \5854 );
mbuf \mul_7_15_g34900/U$1 ( \5857 , \5668 );
mand \mul_7_15_g34644/U$3 ( \5858 , \5856 , \5857 );
mnor \mul_7_15_g34644/U$1 ( \5859 , \5855 , \5858 );
mnot \fopt36909/U$1 ( \5860 , \5859 );
mnot \fopt36908/U$1 ( \5861 , \5860 );
mnot \mul_7_15_g34348/U$3 ( \5862 , \5861 );
mxor \mul_7_15_g34545/U$1 ( \5863 , \5785 , \5724 );
mnot \mul_7_15_g34639/U$1 ( \5864 , \5837 );
mand \mul_7_15_g34502/U$2 ( \5865 , \5863 , \5864 );
mnot \mul_7_15_g34502/U$4 ( \5866 , \5863 );
mand \mul_7_15_g34502/U$3 ( \5867 , \5866 , \5837 );
mnor \mul_7_15_g34502/U$1 ( \5868 , \5865 , \5867 );
mnot \mul_7_15_g34479/U$1 ( \5869 , \5868 );
mnot \mul_7_15_g34348/U$4 ( \5870 , \5869 );
mor \mul_7_15_g34348/U$2 ( \5871 , \5862 , \5870 );
mnot \mul_7_15_g34365/U$3 ( \5872 , \5860 );
mnot \mul_7_15_g34365/U$4 ( \5873 , \5868 );
mor \mul_7_15_g34365/U$2 ( \5874 , \5872 , \5873 );
mxnor \g36536/U$1 ( \5875 , \5744 , \5732 );
mnot \mul_7_15_g35684/U$3 ( \5876 , \4079 );
mnot \mul_7_15_g35684/U$4 ( \5877 , \4107 );
mor \mul_7_15_g35684/U$2 ( \5878 , \5876 , \5877 );
mnand \mul_7_15_g35813/U$1 ( \5879 , \4110 , \5535 );
mnand \mul_7_15_g35684/U$1 ( \5880 , \5878 , \5879 );
mnot \mul_7_15_g35169/U$3 ( \5881 , \5880 );
mnot \mul_7_15_g35169/U$4 ( \5882 , \4302 );
mor \mul_7_15_g35169/U$2 ( \5883 , \5881 , \5882 );
mnand \mul_7_15_g35420/U$1 ( \5884 , \4133 , \5482 );
mnand \mul_7_15_g35169/U$1 ( \5885 , \5883 , \5884 );
mnot \mul_7_15_g35168/U$1 ( \5886 , \5885 );
mnand \mul_7_15_g34861/U$1 ( \5887 , \5875 , \5886 );
mnor \mul_7_15_g35480/U$1 ( \5888 , \4192 , \5418 );
mnot \mul_7_15_g35286/U$3 ( \5889 , \5266 );
mnot \mul_7_15_g35286/U$4 ( \5890 , \5753 );
mor \mul_7_15_g35286/U$2 ( \5891 , \5889 , \5890 );
mnot \mul_7_15_g35738/U$3 ( \5892 , \4094 );
mnot \mul_7_15_g35738/U$4 ( \5893 , \5274 );
mor \mul_7_15_g35738/U$2 ( \5894 , \5892 , \5893 );
mnand \mul_7_15_g35809/U$1 ( \5895 , \5268 , \4298 );
mnand \mul_7_15_g35738/U$1 ( \5896 , \5894 , \5895 );
mnand \mul_7_15_g35463/U$1 ( \5897 , \5271 , \5896 );
mnand \mul_7_15_g35286/U$1 ( \5898 , \5891 , \5897 );
mxor \mul_7_15_g34822/U$4 ( \5899 , \5888 , \5898 );
mnot \g37157/U$3 ( \5900 , \4948 );
mnot \g37157/U$4 ( \5901 , \5737 );
mor \g37157/U$2 ( \5902 , \5900 , \5901 );
mnot \mul_7_15_g35992/U$1 ( \5903 , \2945 );
mand \mul_7_15_g35707/U$2 ( \5904 , \5903 , \4097 );
mnot \mul_7_15_g35972/U$1 ( \5905 , \4853 );
mand \mul_7_15_g35707/U$3 ( \5906 , \5905 , \4254 );
mnor \mul_7_15_g35707/U$1 ( \5907 , \5904 , \5906 );
mnot \g37158/U$2 ( \5908 , \5907 );
mnand \g37158/U$1 ( \5909 , \5908 , \4944 );
mnand \g37157/U$1 ( \5910 , \5902 , \5909 );
mand \mul_7_15_g34822/U$3 ( \5911 , \5899 , \5910 );
mand \mul_7_15_g34822/U$5 ( \5912 , \5888 , \5898 );
mor \mul_7_15_g34822/U$2 ( \5913 , \5911 , \5912 );
mand \mul_7_15_g34728/U$2 ( \5914 , \5887 , \5913 );
mnor \mul_7_15_g34860/U$1 ( \5915 , \5875 , \5886 );
mnor \mul_7_15_g34728/U$1 ( \5916 , \5914 , \5915 );
mnot \mul_7_15_g34638/U$1 ( \5917 , \5916 );
mnot \mul_7_15_g34408/U$3 ( \5918 , \5917 );
mnot \mul_7_15_g35145/U$3 ( \5919 , \4610 );
mnot \mul_7_15_g35656/U$3 ( \5920 , \4095 );
mnot \mul_7_15_g35656/U$4 ( \5921 , \5138 );
mor \mul_7_15_g35656/U$2 ( \5922 , \5920 , \5921 );
mnand \mul_7_15_g35877/U$1 ( \5923 , \4745 , \4391 );
mnand \mul_7_15_g35656/U$1 ( \5924 , \5922 , \5923 );
mnot \mul_7_15_g35145/U$4 ( \5925 , \5924 );
mor \mul_7_15_g35145/U$2 ( \5926 , \5919 , \5925 );
mnand \mul_7_15_g35384/U$1 ( \5927 , \5795 , \5146 );
mnand \mul_7_15_g35145/U$1 ( \5928 , \5926 , \5927 );
mnot \mul_7_15_g34914/U$3 ( \5929 , \5928 );
mnot \mul_7_15_g35153/U$3 ( \5930 , \4450 );
mand \mul_7_15_g35713/U$2 ( \5931 , \4662 , \4458 );
mnot \mul_7_15_g35713/U$4 ( \5932 , \4662 );
mand \mul_7_15_g35713/U$3 ( \5933 , \5932 , \4535 );
mnor \mul_7_15_g35713/U$1 ( \5934 , \5931 , \5933 );
mnot \mul_7_15_g35153/U$4 ( \5935 , \5934 );
mand \mul_7_15_g35153/U$2 ( \5936 , \5930 , \5935 );
mnot \mul_7_15_g36426/U$2 ( \5937 , \4452 );
mnor \mul_7_15_g36426/U$1 ( \5938 , \5937 , \5773 );
mnor \mul_7_15_g35153/U$1 ( \5939 , \5936 , \5938 );
mnot \mul_7_15_g35152/U$1 ( \5940 , \5939 );
mnot \mul_7_15_g34914/U$4 ( \5941 , \5940 );
mor \mul_7_15_g34914/U$2 ( \5942 , \5929 , \5941 );
mnot \mul_7_15_g35144/U$1 ( \5943 , \5928 );
mnot \mul_7_15_g34935/U$3 ( \5944 , \5943 );
mnot \mul_7_15_g34935/U$4 ( \5945 , \5939 );
mor \mul_7_15_g34935/U$2 ( \5946 , \5944 , \5945 );
mnot \mul_7_15_g35669/U$3 ( \5947 , \4026 );
mnot \mul_7_15_g35669/U$4 ( \5948 , \4332 );
mor \mul_7_15_g35669/U$2 ( \5949 , \5947 , \5948 );
mnand \mul_7_15_g35808/U$1 ( \5950 , \4673 , \4969 );
mnand \mul_7_15_g35669/U$1 ( \5951 , \5949 , \5950 );
mnot \mul_7_15_g35159/U$3 ( \5952 , \5951 );
mnot \mul_7_15_g35159/U$4 ( \5953 , \5497 );
mor \mul_7_15_g35159/U$2 ( \5954 , \5952 , \5953 );
mnot \mul_7_15_g36428/U$2 ( \5955 , \5822 );
mnand \mul_7_15_g36428/U$1 ( \5956 , \5955 , \4800 );
mnand \mul_7_15_g35159/U$1 ( \5957 , \5954 , \5956 );
mnand \mul_7_15_g34935/U$1 ( \5958 , \5946 , \5957 );
mnand \mul_7_15_g34914/U$1 ( \5959 , \5942 , \5958 );
mnot \mul_7_15_g34803/U$1 ( \5960 , \5959 );
mnot \fopt36704/U$1 ( \5961 , \5800 );
mnot \mul_7_15_g34974/U$3 ( \5962 , \5961 );
mnot \mul_7_15_g34974/U$4 ( \5963 , \5827 );
mor \mul_7_15_g34974/U$2 ( \5964 , \5962 , \5963 );
mnand \mul_7_15_g34989/U$1 ( \5965 , \5826 , \5800 );
mnand \mul_7_15_g34974/U$1 ( \5966 , \5964 , \5965 );
mand \mul_7_15_g34897/U$2 ( \5967 , \5966 , \5813 );
mnot \mul_7_15_g34897/U$4 ( \5968 , \5966 );
mand \mul_7_15_g34897/U$3 ( \5969 , \5968 , \5814 );
mnor \mul_7_15_g34897/U$1 ( \5970 , \5967 , \5969 );
mnand \mul_7_15_g34736/U$1 ( \5971 , \5960 , \5970 );
mor \mul_7_15_g35025/U$2 ( \5972 , \5907 , \4862 );
mnot \mul_7_15_g35672/U$3 ( \5973 , \4093 );
mnot \mul_7_15_g35971/U$1 ( \5974 , \5905 );
mnot \mul_7_15_g35672/U$4 ( \5975 , \5974 );
mor \mul_7_15_g35672/U$2 ( \5976 , \5973 , \5975 );
mnand \mul_7_15_g35850/U$1 ( \5977 , \5905 , \4349 );
mnand \mul_7_15_g35672/U$1 ( \5978 , \5976 , \5977 );
mnand \mul_7_15_g35267/U$1 ( \5979 , \4862 , \5978 , \4858 );
mnand \mul_7_15_g35025/U$1 ( \5980 , \5972 , \5979 );
mnand \mul_7_15_g35753/U$1 ( \5981 , \4116 , \5418 );
mand \mul_7_15_g35500/U$2 ( \5982 , \4170 , \5981 );
mnot \mul_7_15_g35527/U$3 ( \5983 , \4098 );
mnot \mul_7_15_g35527/U$4 ( \5984 , \4115 );
mor \mul_7_15_g35527/U$2 ( \5985 , \5983 , \5984 );
mnand \mul_7_15_g35527/U$1 ( \5986 , \5985 , \4106 );
mnor \mul_7_15_g35500/U$1 ( \5987 , \5982 , \5986 );
mnand \mul_7_15_g35001/U$1 ( \5988 , \5980 , \5987 );
mnot \mul_7_15_g34723/U$3 ( \5989 , \5988 );
mnot \mul_7_15_g35704/U$3 ( \5990 , \4082 );
mnot \mul_7_15_g35704/U$4 ( \5991 , \4107 );
mor \mul_7_15_g35704/U$2 ( \5992 , \5990 , \5991 );
mnand \mul_7_15_g35838/U$1 ( \5993 , \4110 , \5526 );
mnand \mul_7_15_g35704/U$1 ( \5994 , \5992 , \5993 );
mnot \mul_7_15_g35165/U$3 ( \5995 , \5994 );
mnot \mul_7_15_g35165/U$4 ( \5996 , \4128 );
mor \mul_7_15_g35165/U$2 ( \5997 , \5995 , \5996 );
mnand \mul_7_15_g35349/U$1 ( \5998 , \5880 , \4132 );
mnand \mul_7_15_g35165/U$1 ( \5999 , \5997 , \5998 );
mnot \mul_7_15_g35163/U$1 ( \6000 , \5999 );
mnot \mul_7_15_g34723/U$4 ( \6001 , \6000 );
mor \mul_7_15_g34723/U$2 ( \6002 , \5989 , \6001 );
mnot \mul_7_15_g35637/U$3 ( \6003 , \4076 );
mnot \mul_7_15_g35637/U$4 ( \6004 , \4163 );
mor \mul_7_15_g35637/U$2 ( \6005 , \6003 , \6004 );
mnand \mul_7_15_g35841/U$1 ( \6006 , \4311 , \5284 );
mnand \mul_7_15_g35637/U$1 ( \6007 , \6005 , \6006 );
mnot \mul_7_15_g35161/U$3 ( \6008 , \6007 );
mnot \mul_7_15_g35161/U$4 ( \6009 , \4159 );
mor \mul_7_15_g35161/U$2 ( \6010 , \6008 , \6009 );
mnot \mul_7_15_g36429/U$2 ( \6011 , \5808 );
mnand \mul_7_15_g36429/U$1 ( \6012 , \6011 , \4317 );
mnand \mul_7_15_g35161/U$1 ( \6013 , \6010 , \6012 );
mnand \mul_7_15_g34723/U$1 ( \6014 , \6002 , \6013 );
mnot \mul_7_15_g36396/U$2 ( \6015 , \5988 );
mnand \mul_7_15_g36396/U$1 ( \6016 , \6015 , \5999 );
mnand \mul_7_15_g34685/U$1 ( \6017 , \6014 , \6016 );
mand \mul_7_15_g34582/U$2 ( \6018 , \5971 , \6017 );
mnor \mul_7_15_g34733/U$1 ( \6019 , \5970 , \5960 );
mnor \mul_7_15_g34582/U$1 ( \6020 , \6018 , \6019 );
mnot \mul_7_15_g34516/U$1 ( \6021 , \6020 );
mnot \mul_7_15_g34408/U$4 ( \6022 , \6021 );
mor \mul_7_15_g34408/U$2 ( \6023 , \5918 , \6022 );
mnot \mul_7_15_g34428/U$3 ( \6024 , \5916 );
mnot \mul_7_15_g34428/U$4 ( \6025 , \6020 );
mor \mul_7_15_g34428/U$2 ( \6026 , \6024 , \6025 );
mxor \mul_7_15_g34643/U$1 ( \6027 , \5745 , \5747 );
mxor \mul_7_15_g34643/U$1_r1 ( \6028 , \6027 , \5782 );
mnand \mul_7_15_g34428/U$1 ( \6029 , \6026 , \6028 );
mnand \mul_7_15_g34408/U$1 ( \6030 , \6023 , \6029 );
mnand \mul_7_15_g34365/U$1 ( \6031 , \5874 , \6030 );
mnand \mul_7_15_g34348/U$1 ( \6032 , \5871 , \6031 );
mnor \mul_7_15_g34238/U$1 ( \6033 , \5849 , \6032 );
mnot \fopt36860/U$1 ( \6034 , \6033 );
mnot \mul_7_15_g34303/U$3 ( \6035 , \5868 );
mand \mul_7_15_g36361/U$2 ( \6036 , \5859 , \6030 );
mnot \mul_7_15_g36361/U$4 ( \6037 , \5859 );
mnot \fopt36807/U$1 ( \6038 , \6030 );
mand \mul_7_15_g36361/U$3 ( \6039 , \6037 , \6038 );
mnor \mul_7_15_g36361/U$1 ( \6040 , \6036 , \6039 );
mnot \mul_7_15_g34303/U$4 ( \6041 , \6040 );
mor \mul_7_15_g34303/U$2 ( \6042 , \6035 , \6041 );
mor \mul_7_15_g34303/U$5 ( \6043 , \5868 , \6040 );
mnand \mul_7_15_g34303/U$1 ( \6044 , \6042 , \6043 );
mnot \mul_7_15_g34276/U$1 ( \6045 , \6044 );
mxor \mul_7_15_g34676/U$1 ( \6046 , \5829 , \5834 );
mxnor \mul_7_15_g34676/U$1_r1 ( \6047 , \6046 , \5789 );
mxor \mul_7_15_g34767/U$1 ( \6048 , \5758 , \5768 );
mxor \mul_7_15_g34767/U$1_r1 ( \6049 , \6048 , \5779 );
mxor \mul_7_15_g34822/U$1 ( \6050 , \5888 , \5898 );
mxor \mul_7_15_g34822/U$1_r1 ( \6051 , \6050 , \5910 );
mnot \mul_7_15_g34580/U$3 ( \6052 , \6051 );
mnot \mul_7_15_g35288/U$3 ( \6053 , \5271 );
mnot \mul_7_15_g35735/U$3 ( \6054 , \4096 );
mnot \mul_7_15_g35735/U$4 ( \6055 , \5422 );
mor \mul_7_15_g35735/U$2 ( \6056 , \6054 , \6055 );
mnand \mul_7_15_g35835/U$1 ( \6057 , \4372 , \5268 );
mnand \mul_7_15_g35735/U$1 ( \6058 , \6056 , \6057 );
mnot \mul_7_15_g35288/U$4 ( \6059 , \6058 );
mor \mul_7_15_g35288/U$2 ( \6060 , \6053 , \6059 );
mnand \mul_7_15_g35304/U$1 ( \6061 , \5896 , \5266 );
mnand \mul_7_15_g35288/U$1 ( \6062 , \6060 , \6061 );
mnot \mul_7_15_g34781/U$3 ( \6063 , \6062 );
mnot \mul_7_15_g35134/U$3 ( \6064 , \4449 );
mnot \mul_7_15_g35652/U$3 ( \6065 , \4021 );
mnot \mul_7_15_g35652/U$4 ( \6066 , \4532 );
mor \mul_7_15_g35652/U$2 ( \6067 , \6065 , \6066 );
mnand \mul_7_15_g35849/U$1 ( \6068 , \4458 , \4780 );
mnand \mul_7_15_g35652/U$1 ( \6069 , \6067 , \6068 );
mnot \mul_7_15_g35134/U$4 ( \6070 , \6069 );
mor \mul_7_15_g35134/U$2 ( \6071 , \6064 , \6070 );
mnot \mul_7_15_g36431/U$2 ( \6072 , \5934 );
mnand \mul_7_15_g36431/U$1 ( \6073 , \6072 , \4452 );
mnand \mul_7_15_g35134/U$1 ( \6074 , \6071 , \6073 );
mnot \mul_7_15_g34781/U$4 ( \6075 , \6074 );
mor \mul_7_15_g34781/U$2 ( \6076 , \6063 , \6075 );
mor \mul_7_15_g34872/U$2 ( \6077 , \6074 , \6062 );
mnot \mul_7_15_g35660/U$3 ( \6078 , \4072 );
mnot \mul_7_15_g35660/U$4 ( \6079 , \4284 );
mor \mul_7_15_g35660/U$2 ( \6080 , \6078 , \6079 );
mnand \mul_7_15_g35811/U$1 ( \6081 , \4283 , \5089 );
mnand \mul_7_15_g35660/U$1 ( \6082 , \6080 , \6081 );
mnot \mul_7_15_g35132/U$3 ( \6083 , \6082 );
mnot \mul_7_15_g35132/U$4 ( \6084 , \4797 );
mor \mul_7_15_g35132/U$2 ( \6085 , \6083 , \6084 );
mnot \mul_7_15_g35325/U$2 ( \6086 , \4267 );
mnand \mul_7_15_g35325/U$1 ( \6087 , \6086 , \5951 );
mnand \mul_7_15_g35132/U$1 ( \6088 , \6085 , \6087 );
mnand \mul_7_15_g34872/U$1 ( \6089 , \6077 , \6088 );
mnand \mul_7_15_g34781/U$1 ( \6090 , \6076 , \6089 );
mnot \mul_7_15_g34580/U$4 ( \6091 , \6090 );
mor \mul_7_15_g34580/U$2 ( \6092 , \6052 , \6091 );
mor \mul_7_15_g34621/U$2 ( \6093 , \6051 , \6090 );
mnot \mul_7_15_g35676/U$3 ( \6094 , \4079 );
mnot \mul_7_15_g35676/U$4 ( \6095 , \4163 );
mor \mul_7_15_g35676/U$2 ( \6096 , \6094 , \6095 );
mnand \mul_7_15_g35797/U$1 ( \6097 , \4170 , \5535 );
mnand \mul_7_15_g35676/U$1 ( \6098 , \6096 , \6097 );
mnot \mul_7_15_g35138/U$3 ( \6099 , \6098 );
mnot \mul_7_15_g35138/U$4 ( \6100 , \4159 );
mor \mul_7_15_g35138/U$2 ( \6101 , \6099 , \6100 );
mnand \mul_7_15_g35375/U$1 ( \6102 , \6007 , \4317 );
mnand \mul_7_15_g35138/U$1 ( \6103 , \6101 , \6102 );
mnot \mul_7_15_g35629/U$3 ( \6104 , \4066 );
mnot \mul_7_15_g35629/U$4 ( \6105 , \5138 );
mor \mul_7_15_g35629/U$2 ( \6106 , \6104 , \6105 );
mnand \mul_7_15_g36926/U$1 ( \6107 , \4616 , \4519 );
mnand \mul_7_15_g35629/U$1 ( \6108 , \6106 , \6107 );
mnot \mul_7_15_g35142/U$3 ( \6109 , \6108 );
mnot \mul_7_15_g35142/U$4 ( \6110 , \4611 );
mor \mul_7_15_g35142/U$2 ( \6111 , \6109 , \6110 );
mnand \mul_7_15_g35376/U$1 ( \6112 , \5924 , \4881 );
mnand \mul_7_15_g35142/U$1 ( \6113 , \6111 , \6112 );
mor \mul_7_15_g34934/U$2 ( \6114 , \6103 , \6113 );
mnot \mul_7_15_g35747/U$3 ( \6115 , \4098 );
mnot \mul_7_15_g35747/U$4 ( \6116 , \4206 );
mor \mul_7_15_g35747/U$2 ( \6117 , \6115 , \6116 );
mnand \mul_7_15_g35904/U$1 ( \6118 , \4110 , \5418 );
mnand \mul_7_15_g35747/U$1 ( \6119 , \6117 , \6118 );
mnot \mul_7_15_g35143/U$3 ( \6120 , \6119 );
mnot \mul_7_15_g35143/U$4 ( \6121 , \4710 );
mor \mul_7_15_g35143/U$2 ( \6122 , \6120 , \6121 );
mnand \mul_7_15_g35378/U$1 ( \6123 , \5994 , \4654 );
mnand \mul_7_15_g35143/U$1 ( \6124 , \6122 , \6123 );
mnand \mul_7_15_g34934/U$1 ( \6125 , \6114 , \6124 );
mnand \mul_7_15_g34987/U$1 ( \6126 , \6103 , \6113 );
mnand \mul_7_15_g34911/U$1 ( \6127 , \6125 , \6126 );
mnand \mul_7_15_g34621/U$1 ( \6128 , \6093 , \6127 );
mnand \mul_7_15_g34580/U$1 ( \6129 , \6092 , \6128 );
mxor \mul_7_15_g34478/U$4 ( \6130 , \6049 , \6129 );
mxor \mul_7_15_g34677/U$1 ( \6131 , \5885 , \5913 );
mxnor \mul_7_15_g34677/U$1_r1 ( \6132 , \6131 , \5875 );
mand \mul_7_15_g34478/U$3 ( \6133 , \6130 , \6132 );
mand \mul_7_15_g34478/U$5 ( \6134 , \6049 , \6129 );
mor \mul_7_15_g34478/U$2 ( \6135 , \6133 , \6134 );
mxor \mul_7_15_g34301/U$4 ( \6136 , \6047 , \6135 );
mnot \mul_7_15_g34481/U$3 ( \6137 , \5916 );
mnot \mul_7_15_g34481/U$4 ( \6138 , \6021 );
mor \mul_7_15_g34481/U$2 ( \6139 , \6137 , \6138 );
mnand \mul_7_15_g34484/U$1 ( \6140 , \6020 , \5917 );
mnand \mul_7_15_g34481/U$1 ( \6141 , \6139 , \6140 );
mand \mul_7_15_g34416/U$2 ( \6142 , \6141 , \6028 );
mnot \mul_7_15_g34416/U$4 ( \6143 , \6141 );
mnot \mul_7_15_g34640/U$1 ( \6144 , \6028 );
mand \mul_7_15_g34416/U$3 ( \6145 , \6143 , \6144 );
mnor \mul_7_15_g34416/U$1 ( \6146 , \6142 , \6145 );
mand \mul_7_15_g34301/U$3 ( \6147 , \6136 , \6146 );
mand \mul_7_15_g34301/U$5 ( \6148 , \6047 , \6135 );
mor \mul_7_15_g34301/U$2 ( \6149 , \6147 , \6148 );
mnot \mul_7_15_g34300/U$1 ( \6150 , \6149 );
mnand \mul_7_15_g34239/U$1 ( \6151 , \6045 , \6150 );
mand \mul_7_15_g34608/U$2 ( \6152 , \6017 , \5959 );
mnot \mul_7_15_g34608/U$4 ( \6153 , \6017 );
mand \mul_7_15_g34608/U$3 ( \6154 , \6153 , \5960 );
mnor \mul_7_15_g34608/U$1 ( \6155 , \6152 , \6154 );
mbuf \mul_7_15_g34842/U$1 ( \6156 , \5970 );
mnot \mul_7_15_g34841/U$1 ( \6157 , \6156 );
mand \mul_7_15_g34551/U$2 ( \6158 , \6155 , \6157 );
mnot \mul_7_15_g34551/U$4 ( \6159 , \6155 );
mand \mul_7_15_g34551/U$3 ( \6160 , \6159 , \6156 );
mnor \mul_7_15_g34551/U$1 ( \6161 , \6158 , \6160 );
mxor \g36763/U$1 ( \6162 , \5987 , \5980 );
mnot \mul_7_15_g34737/U$2 ( \6163 , \6162 );
mnot \mul_7_15_g35729/U$3 ( \6164 , \4097 );
mnot \mul_7_15_g35729/U$4 ( \6165 , \5422 );
mor \mul_7_15_g35729/U$2 ( \6166 , \6164 , \6165 );
mnand \mul_7_15_g35890/U$1 ( \6167 , \5268 , \4254 );
mnand \mul_7_15_g35729/U$1 ( \6168 , \6166 , \6167 );
mnot \mul_7_15_g35282/U$3 ( \6169 , \6168 );
mnot \mul_7_15_g35282/U$4 ( \6170 , \5270 );
mor \mul_7_15_g35282/U$2 ( \6171 , \6169 , \6170 );
mnand \mul_7_15_g35365/U$1 ( \6172 , \6058 , \5266 );
mnand \mul_7_15_g35282/U$1 ( \6173 , \6171 , \6172 );
mnot \g37156/U$2 ( \6174 , \6173 );
mnand \mul_7_15_g35475/U$1 ( \6175 , \4132 , \4098 );
mnand \g37156/U$1 ( \6176 , \6174 , \6175 );
mnot \g37155/U$3 ( \6177 , \6176 );
mand \mul_7_15_g35678/U$2 ( \6178 , \4866 , \4095 );
mand \mul_7_15_g35678/U$3 ( \6179 , \4934 , \4391 );
mnor \mul_7_15_g35678/U$1 ( \6180 , \6178 , \6179 );
mnot \mul_7_15_g35677/U$1 ( \6181 , \6180 );
mnot \mul_7_15_g35036/U$3 ( \6182 , \6181 );
mnot \mul_7_15_g35036/U$4 ( \6183 , \4944 );
mor \mul_7_15_g35036/U$2 ( \6184 , \6182 , \6183 );
mnand \mul_7_15_g35379/U$1 ( \6185 , \4863 , \5978 );
mnand \mul_7_15_g35036/U$1 ( \6186 , \6184 , \6185 );
mnot \g37155/U$4 ( \6187 , \6186 );
mor \g37155/U$2 ( \6188 , \6177 , \6187 );
mnot \mul_7_15_g36422/U$2 ( \6189 , \6175 );
mnand \mul_7_15_g36422/U$1 ( \6190 , \6189 , \6173 );
mnand \g37155/U$1 ( \6191 , \6188 , \6190 );
mnot \mul_7_15_g34849/U$1 ( \6192 , \6191 );
mnand \mul_7_15_g34737/U$1 ( \6193 , \6163 , \6192 );
mnot \mul_7_15_g34626/U$3 ( \6194 , \6193 );
mnot \mul_7_15_g35118/U$3 ( \6195 , \4449 );
mnot \mul_7_15_g35638/U$3 ( \6196 , \4026 );
mnot \mul_7_15_g35638/U$4 ( \6197 , \5112 );
mor \mul_7_15_g35638/U$2 ( \6198 , \6196 , \6197 );
mnand \mul_7_15_g35795/U$1 ( \6199 , \4729 , \4969 );
mnand \mul_7_15_g35638/U$1 ( \6200 , \6198 , \6199 );
mnot \mul_7_15_g35118/U$4 ( \6201 , \6200 );
mor \mul_7_15_g35118/U$2 ( \6202 , \6195 , \6201 );
mnand \mul_7_15_g35361/U$1 ( \6203 , \4452 , \6069 );
mnand \mul_7_15_g35118/U$1 ( \6204 , \6202 , \6203 );
mnot \mul_7_15_g35117/U$1 ( \6205 , \6204 );
mnot \mul_7_15_g34933/U$3 ( \6206 , \6205 );
mnot \mul_7_15_g35683/U$3 ( \6207 , \4082 );
mnot \mul_7_15_g35683/U$4 ( \6208 , \4163 );
mor \mul_7_15_g35683/U$2 ( \6209 , \6207 , \6208 );
mnand \mul_7_15_g35857/U$1 ( \6210 , \4170 , \5526 );
mnand \mul_7_15_g35683/U$1 ( \6211 , \6209 , \6210 );
mnot \mul_7_15_g35116/U$3 ( \6212 , \6211 );
mnot \mul_7_15_g35116/U$4 ( \6213 , \4159 );
mor \mul_7_15_g35116/U$2 ( \6214 , \6212 , \6213 );
mnand \mul_7_15_g35360/U$1 ( \6215 , \4317 , \6098 );
mnand \mul_7_15_g35116/U$1 ( \6216 , \6214 , \6215 );
mnot \mul_7_15_g35114/U$1 ( \6217 , \6216 );
mnot \mul_7_15_g34933/U$4 ( \6218 , \6217 );
mor \mul_7_15_g34933/U$2 ( \6219 , \6206 , \6218 );
mnot \mul_7_15_g35634/U$3 ( \6220 , \4076 );
mnot \mul_7_15_g35634/U$4 ( \6221 , \4493 );
mor \mul_7_15_g35634/U$2 ( \6222 , \6220 , \6221 );
mnand \mul_7_15_g35817/U$1 ( \6223 , \4283 , \5284 );
mnand \mul_7_15_g35634/U$1 ( \6224 , \6222 , \6223 );
mnot \mul_7_15_g35120/U$3 ( \6225 , \6224 );
mnot \mul_7_15_g35120/U$4 ( \6226 , \4797 );
mor \mul_7_15_g35120/U$2 ( \6227 , \6225 , \6226 );
mnand \mul_7_15_g35362/U$1 ( \6228 , \6082 , \4800 );
mnand \mul_7_15_g35120/U$1 ( \6229 , \6227 , \6228 );
mnand \mul_7_15_g34933/U$1 ( \6230 , \6219 , \6229 );
mnand \mul_7_15_g34983/U$1 ( \6231 , \6204 , \6216 );
mnand \mul_7_15_g34910/U$1 ( \6232 , \6230 , \6231 );
mnot \mul_7_15_g34626/U$4 ( \6233 , \6232 );
mor \mul_7_15_g34626/U$2 ( \6234 , \6194 , \6233 );
mnand \mul_7_15_g34743/U$1 ( \6235 , \6191 , \6162 );
mnand \mul_7_15_g34626/U$1 ( \6236 , \6234 , \6235 );
mnot \mul_7_15_g34513/U$3 ( \6237 , \6236 );
mnot \mul_7_15_g35151/U$1 ( \6238 , \5940 );
mnot \mul_7_15_g34896/U$3 ( \6239 , \6238 );
mnot \mul_7_15_g34972/U$3 ( \6240 , \5928 );
mnot \mul_7_15_g35158/U$1 ( \6241 , \5957 );
mnot \mul_7_15_g34972/U$4 ( \6242 , \6241 );
mor \mul_7_15_g34972/U$2 ( \6243 , \6240 , \6242 );
mor \mul_7_15_g34972/U$5 ( \6244 , \5928 , \6241 );
mnand \mul_7_15_g34972/U$1 ( \6245 , \6243 , \6244 );
mnot \mul_7_15_g34896/U$4 ( \6246 , \6245 );
mor \mul_7_15_g34896/U$2 ( \6247 , \6239 , \6246 );
mnot \mul_7_15_g34971/U$1 ( \6248 , \6245 );
mnot \mul_7_15_g35150/U$1 ( \6249 , \6238 );
mnand \mul_7_15_g34903/U$1 ( \6250 , \6248 , \6249 );
mnand \mul_7_15_g34896/U$1 ( \6251 , \6247 , \6250 );
mnot \mul_7_15_g36387/U$2 ( \6252 , \6251 );
mand \g37273/U$2 ( \6253 , \5988 , \5999 );
mnot \g37273/U$4 ( \6254 , \5988 );
mand \g37273/U$3 ( \6255 , \6254 , \6000 );
mor \g37273/U$1 ( \6256 , \6253 , \6255 );
mnot \mul_7_15_g35160/U$1 ( \6257 , \6013 );
mand \mul_7_15_g34695/U$2 ( \6258 , \6256 , \6257 );
mnot \mul_7_15_g34695/U$4 ( \6259 , \6256 );
mand \mul_7_15_g34695/U$3 ( \6260 , \6259 , \6013 );
mnor \mul_7_15_g34695/U$1 ( \6261 , \6258 , \6260 );
mnand \mul_7_15_g36387/U$1 ( \6262 , \6252 , \6261 );
mnot \mul_7_15_g34513/U$4 ( \6263 , \6262 );
mor \mul_7_15_g34513/U$2 ( \6264 , \6237 , \6263 );
mnot \mul_7_15_g36374/U$2 ( \6265 , \6261 );
mnand \mul_7_15_g36374/U$1 ( \6266 , \6265 , \6251 );
mnand \mul_7_15_g34513/U$1 ( \6267 , \6264 , \6266 );
mxor \mul_7_15_g34374/U$4 ( \6268 , \6161 , \6267 );
mxor \mul_7_15_g34478/U$1 ( \6269 , \6049 , \6129 );
mxor \mul_7_15_g34478/U$1_r1 ( \6270 , \6269 , \6132 );
mand \mul_7_15_g34374/U$3 ( \6271 , \6268 , \6270 );
mand \mul_7_15_g34374/U$5 ( \6272 , \6161 , \6267 );
mor \mul_7_15_g34374/U$2 ( \6273 , \6271 , \6272 );
mnot \mul_7_15_g34256/U$2 ( \6274 , \6273 );
mxor \mul_7_15_g34301/U$1 ( \6275 , \6047 , \6135 );
mxor \mul_7_15_g34301/U$1_r1 ( \6276 , \6275 , \6146 );
mnot \mul_7_15_g34299/U$1 ( \6277 , \6276 );
mnand \mul_7_15_g34256/U$1 ( \6278 , \6274 , \6277 );
mand \mul_7_15_g34224/U$1 ( \6279 , \6151 , \6278 );
mxor \mul_7_15_g34373/U$1 ( \6280 , \5653 , \5691 );
mxor \mul_7_15_g34373/U$1_r1 ( \6281 , \6280 , \5702 );
mnot \mul_7_15_g34543/U$1 ( \6282 , \5721 );
mnand \mul_7_15_g34437/U$1 ( \6283 , \5847 , \6282 );
mnot \mul_7_15_g34480/U$1 ( \6284 , \5840 );
mand \mul_7_15_g34409/U$2 ( \6285 , \6283 , \6284 );
mnor \mul_7_15_g34436/U$1 ( \6286 , \5847 , \6282 );
mnor \mul_7_15_g34409/U$1 ( \6287 , \6285 , \6286 );
mnand \mul_7_15_g34323/U$1 ( \6288 , \6281 , \6287 );
mnand \mul_7_15_g34218/U$1 ( \6289 , \6034 , \6279 , \6288 );
mnot \mul_7_15_g34217/U$1 ( \6290 , \6289 );
mnot \mul_7_15_g35691/U$3 ( \6291 , \4082 );
mnot \mul_7_15_g35691/U$4 ( \6292 , \5301 );
mor \mul_7_15_g35691/U$2 ( \6293 , \6291 , \6292 );
mnand \mul_7_15_g35873/U$1 ( \6294 , \4616 , \5526 );
mnand \mul_7_15_g35691/U$1 ( \6295 , \6293 , \6294 );
mnot \mul_7_15_g35079/U$3 ( \6296 , \6295 );
mnot \mul_7_15_g35079/U$4 ( \6297 , \4611 );
mor \mul_7_15_g35079/U$2 ( \6298 , \6296 , \6297 );
mnot \mul_7_15_g35682/U$3 ( \6299 , \4079 );
mnot \mul_7_15_g35682/U$4 ( \6300 , \5301 );
mor \mul_7_15_g35682/U$2 ( \6301 , \6299 , \6300 );
mnot \mul_7_15_g36436/U$2 ( \6302 , \5138 );
mnand \mul_7_15_g36436/U$1 ( \6303 , \6302 , \5535 );
mnand \mul_7_15_g35682/U$1 ( \6304 , \6301 , \6303 );
mnand \mul_7_15_g35380/U$1 ( \6305 , \6304 , \5146 );
mnand \mul_7_15_g35079/U$1 ( \6306 , \6298 , \6305 );
mnot \mul_7_15_g36402/U$2 ( \6307 , \6306 );
mnot \mul_7_15_g35688/U$3 ( \6308 , \4079 );
mnot \mul_7_15_g35688/U$4 ( \6309 , \4939 );
mor \mul_7_15_g35688/U$2 ( \6310 , \6308 , \6309 );
mnand \mul_7_15_g35794/U$1 ( \6311 , \4936 , \5535 );
mnand \mul_7_15_g35688/U$1 ( \6312 , \6310 , \6311 );
mnot \mul_7_15_g35040/U$3 ( \6313 , \6312 );
mnot \mul_7_15_g35040/U$4 ( \6314 , \4945 );
mor \mul_7_15_g35040/U$2 ( \6315 , \6313 , \6314 );
mand \mul_7_15_g35705/U$2 ( \6316 , \4076 , \4949 );
mnot \mul_7_15_g35705/U$4 ( \6317 , \4076 );
mand \mul_7_15_g35705/U$3 ( \6318 , \6317 , \4935 );
mnor \mul_7_15_g35705/U$1 ( \6319 , \6316 , \6318 );
mnand \mul_7_15_g35404/U$1 ( \6320 , \4948 , \6319 );
mnand \mul_7_15_g35040/U$1 ( \6321 , \6315 , \6320 );
mnot \mul_7_15_g35524/U$3 ( \6322 , \5418 );
mnot \mul_7_15_g35524/U$4 ( \6323 , \4597 );
mor \mul_7_15_g35524/U$2 ( \6324 , \6322 , \6323 );
mnand \mul_7_15_g35524/U$1 ( \6325 , \6324 , \4868 );
mnand \mul_7_15_g35758/U$1 ( \6326 , \3516 , \4098 );
mand \mul_7_15_g35505/U$1 ( \6327 , \6325 , \4616 , \6326 );
mnand \mul_7_15_g35002/U$1 ( \6328 , \6321 , \6327 );
mnand \mul_7_15_g36402/U$1 ( \6329 , \6307 , \6328 );
mnot \mul_7_15_g34682/U$3 ( \6330 , \6329 );
mnot \mul_7_15_g35742/U$3 ( \6331 , \4026 );
mnot \mul_7_15_g35742/U$4 ( \6332 , \5274 );
mor \mul_7_15_g35742/U$2 ( \6333 , \6331 , \6332 );
mnand \mul_7_15_g35881/U$1 ( \6334 , \5425 , \4969 );
mnand \mul_7_15_g35742/U$1 ( \6335 , \6333 , \6334 );
mnot \mul_7_15_g35290/U$3 ( \6336 , \6335 );
mnot \mul_7_15_g35895/U$1 ( \6337 , \5272 );
mnot \mul_7_15_g35290/U$4 ( \6338 , \6337 );
mor \mul_7_15_g35290/U$2 ( \6339 , \6336 , \6338 );
mnot \mul_7_15_g35739/U$3 ( \6340 , \4021 );
mnot \mul_7_15_g35739/U$4 ( \6341 , \5274 );
mor \mul_7_15_g35739/U$2 ( \6342 , \6340 , \6341 );
mnand \mul_7_15_g35820/U$1 ( \6343 , \5425 , \4780 );
mnand \mul_7_15_g35739/U$1 ( \6344 , \6342 , \6343 );
mnand \mul_7_15_g35317/U$1 ( \6345 , \6344 , \5266 );
mnand \mul_7_15_g35290/U$1 ( \6346 , \6339 , \6345 );
mnor \mul_7_15_g35481/U$1 ( \6347 , \4454 , \5418 );
mxor \mul_7_15_g34827/U$1 ( \6348 , \6346 , \6347 );
mnot \mul_7_15_g35035/U$3 ( \6349 , \4945 );
mnot \mul_7_15_g35035/U$4 ( \6350 , \6319 );
mor \mul_7_15_g35035/U$2 ( \6351 , \6349 , \6350 );
mnot \mul_7_15_g35653/U$3 ( \6352 , \4072 );
mnot \mul_7_15_g35653/U$4 ( \6353 , \4869 );
mor \mul_7_15_g35653/U$2 ( \6354 , \6352 , \6353 );
mnand \mul_7_15_g35869/U$1 ( \6355 , \4868 , \5089 );
mnand \mul_7_15_g35653/U$1 ( \6356 , \6354 , \6355 );
mnand \mul_7_15_g35340/U$1 ( \6357 , \4948 , \6356 );
mnand \mul_7_15_g35035/U$1 ( \6358 , \6351 , \6357 );
mxor \mul_7_15_g34827/U$1_r1 ( \6359 , \6348 , \6358 );
mnot \mul_7_15_g34682/U$4 ( \6360 , \6359 );
mor \mul_7_15_g34682/U$2 ( \6361 , \6330 , \6360 );
mnot \mul_7_15_g36395/U$2 ( \6362 , \6328 );
mnand \mul_7_15_g36395/U$1 ( \6363 , \6362 , \6306 );
mnand \mul_7_15_g34682/U$1 ( \6364 , \6361 , \6363 );
mnand \mul_7_15_g35755/U$1 ( \6365 , \4437 , \5418 );
mand \mul_7_15_g35502/U$2 ( \6366 , \4616 , \6365 );
mnot \mul_7_15_g35526/U$3 ( \6367 , \4098 );
mnot \mul_7_15_g36013/U$1 ( \6368 , \4437 );
mnot \mul_7_15_g35526/U$4 ( \6369 , \6368 );
mor \mul_7_15_g35526/U$2 ( \6370 , \6367 , \6369 );
mnand \mul_7_15_g35526/U$1 ( \6371 , \6370 , \4729 );
mnor \mul_7_15_g35502/U$1 ( \6372 , \6366 , \6371 );
mnot \mul_7_15_g35501/U$1 ( \6373 , \6372 );
mnot \mul_7_15_g34960/U$3 ( \6374 , \6373 );
mnot \mul_7_15_g35047/U$3 ( \6375 , \6356 );
mnot \mul_7_15_g35047/U$4 ( \6376 , \4945 );
mor \mul_7_15_g35047/U$2 ( \6377 , \6375 , \6376 );
mnot \mul_7_15_g35680/U$3 ( \6378 , \4026 );
mnot \mul_7_15_g35680/U$4 ( \6379 , \4935 );
mor \mul_7_15_g35680/U$2 ( \6380 , \6378 , \6379 );
mnand \mul_7_15_g35880/U$1 ( \6381 , \2945 , \4969 );
mnand \mul_7_15_g35680/U$1 ( \6382 , \6380 , \6381 );
mnand \mul_7_15_g35389/U$1 ( \6383 , \4863 , \6382 );
mnand \mul_7_15_g35047/U$1 ( \6384 , \6377 , \6383 );
mnot \mul_7_15_g34960/U$4 ( \6385 , \6384 );
mor \mul_7_15_g34960/U$2 ( \6386 , \6374 , \6385 );
mor \mul_7_15_g34960/U$5 ( \6387 , \6384 , \6373 );
mnand \mul_7_15_g34960/U$1 ( \6388 , \6386 , \6387 );
mxor \mul_7_15_g34827/U$4 ( \6389 , \6346 , \6347 );
mand \mul_7_15_g34827/U$3 ( \6390 , \6389 , \6358 );
mand \mul_7_15_g34827/U$5 ( \6391 , \6346 , \6347 );
mor \mul_7_15_g34827/U$2 ( \6392 , \6390 , \6391 );
mxor \mul_7_15_g34594/U$1 ( \6393 , \6388 , \6392 );
mnot \mul_7_15_g35299/U$3 ( \6394 , \6344 );
mnot \mul_7_15_g35299/U$4 ( \6395 , \6337 );
mor \mul_7_15_g35299/U$2 ( \6396 , \6394 , \6395 );
mnot \mul_7_15_g35732/U$3 ( \6397 , \4017 );
mnot \mul_7_15_g35732/U$4 ( \6398 , \5422 );
mor \mul_7_15_g35732/U$2 ( \6399 , \6397 , \6398 );
mnand \mul_7_15_g35831/U$1 ( \6400 , \4662 , \5275 );
mnand \mul_7_15_g35732/U$1 ( \6401 , \6399 , \6400 );
mnand \mul_7_15_g35424/U$1 ( \6402 , \6401 , \5266 );
mnand \mul_7_15_g35299/U$1 ( \6403 , \6396 , \6402 );
mnot \mul_7_15_g35077/U$3 ( \6404 , \6304 );
mnot \mul_7_15_g35077/U$4 ( \6405 , \4611 );
mor \mul_7_15_g35077/U$2 ( \6406 , \6404 , \6405 );
mand \mul_7_15_g35622/U$2 ( \6407 , \4076 , \4616 );
mnot \mul_7_15_g35622/U$4 ( \6408 , \4076 );
mand \mul_7_15_g35622/U$3 ( \6409 , \6408 , \5138 );
mnor \mul_7_15_g35622/U$1 ( \6410 , \6407 , \6409 );
mnand \mul_7_15_g35434/U$1 ( \6411 , \6410 , \4754 );
mnand \mul_7_15_g35077/U$1 ( \6412 , \6406 , \6411 );
mxor \mul_7_15_g34812/U$1 ( \6413 , \6403 , \6412 );
mand \mul_7_15_g35750/U$2 ( \6414 , \4098 , \4532 );
mnot \mul_7_15_g35750/U$4 ( \6415 , \4098 );
mand \mul_7_15_g35750/U$3 ( \6416 , \6415 , \4458 );
mnor \mul_7_15_g35750/U$1 ( \6417 , \6414 , \6416 );
mnot \mul_7_15_g35320/U$1 ( \6418 , \4632 );
mor \mul_7_15_g35179/U$2 ( \6419 , \6417 , \6418 );
mand \mul_7_15_g35686/U$2 ( \6420 , \4082 , \4917 );
mnot \mul_7_15_g35686/U$4 ( \6421 , \4082 );
mand \mul_7_15_g35686/U$3 ( \6422 , \6421 , \4535 );
mnor \mul_7_15_g35686/U$1 ( \6423 , \6420 , \6422 );
mnot \mul_7_15_g35685/U$1 ( \6424 , \6423 );
mor \mul_7_15_g35179/U$3 ( \6425 , \4454 , \6424 );
mnand \mul_7_15_g35179/U$1 ( \6426 , \6419 , \6425 );
mxor \mul_7_15_g34812/U$1_r1 ( \6427 , \6413 , \6426 );
mxor \mul_7_15_g34594/U$1_r1 ( \6428 , \6393 , \6427 );
mxor \mul_7_15_g34389/U$4 ( \6429 , \6364 , \6428 );
mnot \mul_7_15_g35748/U$3 ( \6430 , \5418 );
mnot \mul_7_15_g35748/U$4 ( \6431 , \4616 );
mor \mul_7_15_g35748/U$2 ( \6432 , \6430 , \6431 );
mnand \mul_7_15_g35901/U$1 ( \6433 , \5301 , \4098 );
mnand \mul_7_15_g35748/U$1 ( \6434 , \6432 , \6433 );
mnot \mul_7_15_g35189/U$3 ( \6435 , \6434 );
mnot \mul_7_15_g35189/U$4 ( \6436 , \4611 );
mor \mul_7_15_g35189/U$2 ( \6437 , \6435 , \6436 );
mnand \mul_7_15_g35316/U$1 ( \6438 , \6295 , \4754 );
mnand \mul_7_15_g35189/U$1 ( \6439 , \6437 , \6438 );
mnot \mul_7_15_g36411/U$2 ( \6440 , \6439 );
mnot \mul_7_15_g35736/U$3 ( \6441 , \4072 );
mnot \mul_7_15_g35736/U$4 ( \6442 , \5422 );
mor \mul_7_15_g35736/U$2 ( \6443 , \6441 , \6442 );
mnand \mul_7_15_g35840/U$1 ( \6444 , \5275 , \5089 );
mnand \mul_7_15_g35736/U$1 ( \6445 , \6443 , \6444 );
mnot \mul_7_15_g35295/U$3 ( \6446 , \6445 );
mnot \mul_7_15_g35295/U$4 ( \6447 , \6337 );
mor \mul_7_15_g35295/U$2 ( \6448 , \6446 , \6447 );
mnand \mul_7_15_g35435/U$1 ( \6449 , \6335 , \5266 );
mnand \mul_7_15_g35295/U$1 ( \6450 , \6448 , \6449 );
mnot \mul_7_15_g35294/U$1 ( \6451 , \6450 );
mnand \mul_7_15_g36411/U$1 ( \6452 , \6440 , \6451 );
mnot \mul_7_15_g34782/U$3 ( \6453 , \6452 );
mnot \mul_7_15_g34961/U$3 ( \6454 , \6327 );
mnot \mul_7_15_g35039/U$1 ( \6455 , \6321 );
mnot \mul_7_15_g34961/U$4 ( \6456 , \6455 );
mor \mul_7_15_g34961/U$2 ( \6457 , \6454 , \6456 );
mor \mul_7_15_g34961/U$5 ( \6458 , \6455 , \6327 );
mnand \mul_7_15_g34961/U$1 ( \6459 , \6457 , \6458 );
mnot \mul_7_15_g34782/U$4 ( \6460 , \6459 );
mor \mul_7_15_g34782/U$2 ( \6461 , \6453 , \6460 );
mnand \mul_7_15_g34997/U$1 ( \6462 , \6439 , \6450 );
mnand \mul_7_15_g34782/U$1 ( \6463 , \6461 , \6462 );
mnot \mul_7_15_g36382/U$2 ( \6464 , \6463 );
mnot \mul_7_15_g34791/U$3 ( \6465 , \6328 );
mnot \mul_7_15_g34791/U$4 ( \6466 , \6306 );
mand \mul_7_15_g34791/U$2 ( \6467 , \6465 , \6466 );
mand \mul_7_15_g34791/U$5 ( \6468 , \6328 , \6306 );
mnor \mul_7_15_g34791/U$1 ( \6469 , \6467 , \6468 );
mxor \mul_7_15_g36391/U$1 ( \6470 , \6359 , \6469 );
mnand \mul_7_15_g36382/U$1 ( \6471 , \6464 , \6470 );
mnot \mul_7_15_g34470/U$3 ( \6472 , \6471 );
mnot \mul_7_15_g35477/U$2 ( \6473 , \4602 );
mnand \mul_7_15_g35477/U$1 ( \6474 , \6473 , \4098 );
mnot \mul_7_15_g35726/U$3 ( \6475 , \4082 );
mnot \mul_7_15_g35726/U$4 ( \6476 , \4939 );
mor \mul_7_15_g35726/U$2 ( \6477 , \6475 , \6476 );
mnand \mul_7_15_g35812/U$1 ( \6478 , \4936 , \5526 );
mnand \mul_7_15_g35726/U$1 ( \6479 , \6477 , \6478 );
mnot \mul_7_15_g35048/U$3 ( \6480 , \6479 );
mnot \mul_7_15_g35048/U$4 ( \6481 , \4945 );
mor \mul_7_15_g35048/U$2 ( \6482 , \6480 , \6481 );
mnand \mul_7_15_g35334/U$1 ( \6483 , \6312 , \4863 );
mnand \mul_7_15_g35048/U$1 ( \6484 , \6482 , \6483 );
mxor \mul_7_15_g34887/U$1 ( \6485 , \6474 , \6484 );
mnot \mul_7_15_g35734/U$3 ( \6486 , \4076 );
mnot \mul_7_15_g35734/U$4 ( \6487 , \5422 );
mor \mul_7_15_g35734/U$2 ( \6488 , \6486 , \6487 );
mnand \mul_7_15_g35882/U$1 ( \6489 , \5425 , \5284 );
mnand \mul_7_15_g35734/U$1 ( \6490 , \6488 , \6489 );
mnot \mul_7_15_g35894/U$1 ( \6491 , \5270 );
mnot \mul_7_15_g35892/U$1 ( \6492 , \6491 );
mnand \mul_7_15_g35437/U$1 ( \6493 , \6490 , \6492 );
mnand \mul_7_15_g35355/U$1 ( \6494 , \5266 , \6445 );
mand \mul_7_15_g35277/U$1 ( \6495 , \6493 , \6494 );
mxnor \mul_7_15_g34887/U$1_r1 ( \6496 , \6485 , \6495 );
mnand \mul_7_15_g35756/U$1 ( \6497 , \4851 , \4098 );
mand \mul_7_15_g35525/U$1 ( \6498 , \4934 , \6497 );
mnot \mul_7_15_g35521/U$3 ( \6499 , \5418 );
mnot \mul_7_15_g35521/U$4 ( \6500 , \4856 );
mor \mul_7_15_g35521/U$2 ( \6501 , \6499 , \6500 );
mnand \mul_7_15_g35521/U$1 ( \6502 , \6501 , \5275 );
mnand \mul_7_15_g35504/U$1 ( \6503 , \6498 , \6502 );
mnot \mul_7_15_g36423/U$2 ( \6504 , \6503 );
mand \mul_7_15_g35749/U$2 ( \6505 , \5418 , \4935 );
mnot \mul_7_15_g35749/U$4 ( \6506 , \5418 );
mand \mul_7_15_g35749/U$3 ( \6507 , \6506 , \4949 );
mnor \mul_7_15_g35749/U$1 ( \6508 , \6505 , \6507 );
mnot \mul_7_15_g35050/U$3 ( \6509 , \6508 );
mnot \mul_7_15_g35050/U$4 ( \6510 , \4945 );
mor \mul_7_15_g35050/U$2 ( \6511 , \6509 , \6510 );
mnand \mul_7_15_g35462/U$1 ( \6512 , \4948 , \6479 );
mnand \mul_7_15_g35050/U$1 ( \6513 , \6511 , \6512 );
mnand \mul_7_15_g36423/U$1 ( \6514 , \6504 , \6513 );
mnand \mul_7_15_g34742/U$1 ( \6515 , \6496 , \6514 );
mnot \mul_7_15_g34625/U$3 ( \6516 , \6515 );
mnot \mul_7_15_g35727/U$3 ( \6517 , \5535 );
mnot \mul_7_15_g35727/U$4 ( \6518 , \5275 );
mor \mul_7_15_g35727/U$2 ( \6519 , \6517 , \6518 );
mnand \mul_7_15_g35888/U$1 ( \6520 , \5422 , \4079 );
mnand \mul_7_15_g35727/U$1 ( \6521 , \6519 , \6520 );
mnot \mul_7_15_g35275/U$3 ( \6522 , \6521 );
mnot \mul_7_15_g35275/U$4 ( \6523 , \6337 );
mor \mul_7_15_g35275/U$2 ( \6524 , \6522 , \6523 );
mnand \mul_7_15_g35335/U$1 ( \6525 , \6490 , \5266 );
mnand \mul_7_15_g35275/U$1 ( \6526 , \6524 , \6525 );
mnot \mul_7_15_g35741/U$3 ( \6527 , \4082 );
mnot \mul_7_15_g35741/U$4 ( \6528 , \5274 );
mor \mul_7_15_g35741/U$2 ( \6529 , \6527 , \6528 );
mnand \mul_7_15_g35814/U$1 ( \6530 , \5433 , \5526 );
mnand \mul_7_15_g35741/U$1 ( \6531 , \6529 , \6530 );
mnot \mul_7_15_g35740/U$1 ( \6532 , \6531 );
mnot \mul_7_15_g35301/U$3 ( \6533 , \6532 );
mnot \mul_7_15_g35301/U$4 ( \6534 , \6491 );
mand \mul_7_15_g35301/U$2 ( \6535 , \6533 , \6534 );
mand \mul_7_15_g35301/U$5 ( \6536 , \6521 , \5266 );
mnor \mul_7_15_g35301/U$1 ( \6537 , \6535 , \6536 );
mnand \mul_7_15_g35473/U$1 ( \6538 , \4863 , \4098 );
mnand \mul_7_15_g35016/U$1 ( \6539 , \6537 , \6538 );
mnot \mul_7_15_g35283/U$3 ( \6540 , \5271 );
mnot \mul_7_15_fopt36312/U$1 ( \6541 , \5433 );
mand \mul_7_15_g35751/U$2 ( \6542 , \5418 , \6541 );
mnot \mul_7_15_g35751/U$4 ( \6543 , \5418 );
mand \mul_7_15_g35751/U$3 ( \6544 , \6543 , \5275 );
mnor \mul_7_15_g35751/U$1 ( \6545 , \6542 , \6544 );
mnot \mul_7_15_g35283/U$4 ( \6546 , \6545 );
mor \mul_7_15_g35283/U$2 ( \6547 , \6540 , \6546 );
mnand \mul_7_15_g35461/U$1 ( \6548 , \6531 , \5266 );
mnand \mul_7_15_g35283/U$1 ( \6549 , \6547 , \6548 );
mnand \mul_7_15_g35785/U$1 ( \6550 , \5266 , \4098 );
mand \g37044/U$1 ( \6551 , \6550 , \5425 );
mnand \mul_7_15_g35010/U$1 ( \6552 , \6549 , \6551 );
mnot \mul_7_15_g34963/U$1 ( \6553 , \6552 );
mnand \mul_7_15_g34904/U$1 ( \6554 , \6539 , \6553 );
mnot \mul_7_15_g35300/U$1 ( \6555 , \6537 );
mnot \mul_7_15_g35472/U$1 ( \6556 , \6538 );
mnand \mul_7_15_g35015/U$1 ( \6557 , \6555 , \6556 );
mnand \mul_7_15_g34882/U$1 ( \6558 , \6554 , \6557 );
mxor \mul_7_15_g34698/U$4 ( \6559 , \6526 , \6558 );
mnot \mul_7_15_g34956/U$3 ( \6560 , \6503 );
mnot \mul_7_15_g34956/U$4 ( \6561 , \6513 );
mor \mul_7_15_g34956/U$2 ( \6562 , \6560 , \6561 );
mor \mul_7_15_g34956/U$5 ( \6563 , \6513 , \6503 );
mnand \mul_7_15_g34956/U$1 ( \6564 , \6562 , \6563 );
mand \mul_7_15_g34698/U$3 ( \6565 , \6559 , \6564 );
mand \mul_7_15_g34698/U$5 ( \6566 , \6526 , \6558 );
mor \mul_7_15_g34698/U$2 ( \6567 , \6565 , \6566 );
mnot \mul_7_15_g34625/U$4 ( \6568 , \6567 );
mor \mul_7_15_g34625/U$2 ( \6569 , \6516 , \6568 );
mor \mul_7_15_g36388/U$1 ( \6570 , \6496 , \6514 );
mnand \mul_7_15_g34625/U$1 ( \6571 , \6569 , \6570 );
mnot \mul_7_15_g35006/U$3 ( \6572 , \6474 );
mnot \mul_7_15_g35006/U$4 ( \6573 , \6495 );
mor \mul_7_15_g35006/U$2 ( \6574 , \6572 , \6573 );
mnand \mul_7_15_g35006/U$1 ( \6575 , \6574 , \6484 );
mor \mul_7_15_g36419/U$1 ( \6576 , \6495 , \6474 );
mnand \mul_7_15_g34945/U$1 ( \6577 , \6575 , \6576 );
mnot \mul_7_15_g34711/U$2 ( \6578 , \6577 );
mnot \mul_7_15_g34855/U$3 ( \6579 , \6459 );
mnot \mul_7_15_g34955/U$3 ( \6580 , \6439 );
mnot \mul_7_15_g34955/U$4 ( \6581 , \6451 );
mand \mul_7_15_g34955/U$2 ( \6582 , \6580 , \6581 );
mand \mul_7_15_g34955/U$5 ( \6583 , \6439 , \6451 );
mnor \mul_7_15_g34955/U$1 ( \6584 , \6582 , \6583 );
mnot \mul_7_15_g34855/U$4 ( \6585 , \6584 );
mand \mul_7_15_g34855/U$2 ( \6586 , \6579 , \6585 );
mand \mul_7_15_g34855/U$5 ( \6587 , \6459 , \6584 );
mnor \mul_7_15_g34855/U$1 ( \6588 , \6586 , \6587 );
mnand \mul_7_15_g34711/U$1 ( \6589 , \6578 , \6588 );
mnand \mul_7_15_g34558/U$1 ( \6590 , \6571 , \6589 );
mnot \mul_7_15_g34759/U$1 ( \6591 , \6588 );
mnand \mul_7_15_g34707/U$1 ( \6592 , \6591 , \6577 );
mnand \mul_7_15_g34533/U$1 ( \6593 , \6590 , \6592 );
mnot \mul_7_15_g34470/U$4 ( \6594 , \6593 );
mor \mul_7_15_g34470/U$2 ( \6595 , \6472 , \6594 );
mnot \mul_7_15_g36373/U$2 ( \6596 , \6470 );
mnand \mul_7_15_g36373/U$1 ( \6597 , \6596 , \6463 );
mnand \mul_7_15_g34470/U$1 ( \6598 , \6595 , \6597 );
mand \mul_7_15_g34389/U$3 ( \6599 , \6429 , \6598 );
mand \mul_7_15_g34389/U$5 ( \6600 , \6364 , \6428 );
mor \mul_7_15_g34389/U$2 ( \6601 , \6599 , \6600 );
mnot \mul_7_15_g34344/U$3 ( \6602 , \6601 );
mnot \mul_7_15_g35646/U$3 ( \6603 , \5089 );
mnot \mul_7_15_g35646/U$4 ( \6604 , \4729 );
mor \mul_7_15_g35646/U$2 ( \6605 , \6603 , \6604 );
mnand \mul_7_15_g35823/U$1 ( \6606 , \4457 , \4072 );
mnand \mul_7_15_g35646/U$1 ( \6607 , \6605 , \6606 );
mnot \mul_7_15_g35109/U$3 ( \6608 , \6607 );
mnot \mul_7_15_g35109/U$4 ( \6609 , \4449 );
mor \mul_7_15_g35109/U$2 ( \6610 , \6608 , \6609 );
mnand \mul_7_15_g35342/U$1 ( \6611 , \6200 , \4452 );
mnand \mul_7_15_g35109/U$1 ( \6612 , \6610 , \6611 );
mnot \mul_7_15_g35737/U$3 ( \6613 , \4093 );
mnot \mul_7_15_g35737/U$4 ( \6614 , \5422 );
mor \mul_7_15_g35737/U$2 ( \6615 , \6613 , \6614 );
mnand \mul_7_15_g35816/U$1 ( \6616 , \5433 , \4349 );
mnand \mul_7_15_g35737/U$1 ( \6617 , \6615 , \6616 );
mnot \mul_7_15_g35285/U$3 ( \6618 , \6617 );
mnot \mul_7_15_g35285/U$4 ( \6619 , \6492 );
mor \mul_7_15_g35285/U$2 ( \6620 , \6618 , \6619 );
mnand \mul_7_15_g35347/U$1 ( \6621 , \6168 , \5266 );
mnand \mul_7_15_g35285/U$1 ( \6622 , \6620 , \6621 );
mxor \mul_7_15_g36420/U$1 ( \6623 , \6612 , \6622 );
mnot \mul_7_15_g35642/U$3 ( \6624 , \4079 );
mnot \mul_7_15_g35642/U$4 ( \6625 , \4493 );
mor \mul_7_15_g35642/U$2 ( \6626 , \6624 , \6625 );
mnand \mul_7_15_g35829/U$1 ( \6627 , \4283 , \5535 );
mnand \mul_7_15_g35642/U$1 ( \6628 , \6626 , \6627 );
mnot \mul_7_15_g35105/U$3 ( \6629 , \6628 );
mnot \mul_7_15_g35105/U$4 ( \6630 , \4338 );
mor \mul_7_15_g35105/U$2 ( \6631 , \6629 , \6630 );
mnand \mul_7_15_g35345/U$1 ( \6632 , \5160 , \6224 );
mnand \mul_7_15_g35105/U$1 ( \6633 , \6631 , \6632 );
mxor \mul_7_15_g34853/U$1 ( \6634 , \6623 , \6633 );
mnot \mul_7_15_g34550/U$3 ( \6635 , \6634 );
mnot \mul_7_15_g35024/U$3 ( \6636 , \4862 );
mand \mul_7_15_g35655/U$2 ( \6637 , \4866 , \4017 );
mand \mul_7_15_g35655/U$3 ( \6638 , \4934 , \4662 );
mnor \mul_7_15_g35655/U$1 ( \6639 , \6637 , \6638 );
mnot \mul_7_15_g35024/U$4 ( \6640 , \6639 );
mand \mul_7_15_g35024/U$2 ( \6641 , \6636 , \6640 );
mnot \mul_7_15_g35628/U$3 ( \6642 , \4021 );
mnot \mul_7_15_g35628/U$4 ( \6643 , \4939 );
mor \mul_7_15_g35628/U$2 ( \6644 , \6642 , \6643 );
mnand \mul_7_15_g35862/U$1 ( \6645 , \4867 , \4780 );
mnand \mul_7_15_g35628/U$1 ( \6646 , \6644 , \6645 );
mnand \mul_7_15_g35433/U$1 ( \6647 , \6646 , \4859 );
mnot \mul_7_15_g35432/U$1 ( \6648 , \6647 );
mand \mul_7_15_g35024/U$5 ( \6649 , \6648 , \4862 );
mnor \mul_7_15_g35024/U$1 ( \6650 , \6641 , \6649 );
mnot \mul_7_15_g35523/U$3 ( \6651 , \5418 );
mnot \mul_7_15_g35523/U$4 ( \6652 , \4270 );
mor \mul_7_15_g35523/U$2 ( \6653 , \6651 , \6652 );
mnand \mul_7_15_g35523/U$1 ( \6654 , \6653 , \4917 );
mnand \mul_7_15_g35757/U$1 ( \6655 , \4274 , \4098 );
mnand \mul_7_15_g35496/U$1 ( \6656 , \6654 , \4285 , \6655 );
mor \mul_7_15_g36399/U$1 ( \6657 , \6650 , \6656 );
mnot \mul_7_15_g34651/U$3 ( \6658 , \6657 );
mnand \mul_7_15_g35485/U$1 ( \6659 , \4150 , \4098 );
mnot \mul_7_15_g35484/U$1 ( \6660 , \6659 );
mnot \mul_7_15_g35733/U$3 ( \6661 , \4095 );
mnot \mul_7_15_g35733/U$4 ( \6662 , \5274 );
mor \mul_7_15_g35733/U$2 ( \6663 , \6661 , \6662 );
mnand \mul_7_15_g35859/U$1 ( \6664 , \5433 , \4391 );
mnand \mul_7_15_g35733/U$1 ( \6665 , \6663 , \6664 );
mnot \mul_7_15_g35274/U$3 ( \6666 , \6665 );
mnot \mul_7_15_g35274/U$4 ( \6667 , \5270 );
mor \mul_7_15_g35274/U$2 ( \6668 , \6666 , \6667 );
mnand \mul_7_15_g35430/U$1 ( \6669 , \6617 , \5266 );
mnand \mul_7_15_g35274/U$1 ( \6670 , \6668 , \6669 );
mand \mul_7_15_g3/U$2 ( \6671 , \6660 , \6670 );
mnot \mul_7_15_g3/U$4 ( \6672 , \6660 );
mnot \mul_7_15_g35273/U$1 ( \6673 , \6670 );
mand \mul_7_15_g3/U$3 ( \6674 , \6672 , \6673 );
mnor \mul_7_15_g3/U$1 ( \6675 , \6671 , \6674 );
mnot \mul_7_15_g35654/U$1 ( \6676 , \6639 );
mnot \mul_7_15_g35034/U$3 ( \6677 , \6676 );
mnot \mul_7_15_g35034/U$4 ( \6678 , \4945 );
mor \mul_7_15_g35034/U$2 ( \6679 , \6677 , \6678 );
mnot \mul_7_15_g35658/U$3 ( \6680 , \4066 );
mnot \mul_7_15_g35658/U$4 ( \6681 , \5903 );
mor \mul_7_15_g35658/U$2 ( \6682 , \6680 , \6681 );
mnand \mul_7_15_g35807/U$1 ( \6683 , \5905 , \4519 );
mnand \mul_7_15_g35658/U$1 ( \6684 , \6682 , \6683 );
mnand \mul_7_15_g35328/U$1 ( \6685 , \4948 , \6684 );
mnand \mul_7_15_g35034/U$1 ( \6686 , \6679 , \6685 );
mnot \mul_7_15_g35033/U$1 ( \6687 , \6686 );
mxor \mul_7_15_g36333/U$1 ( \6688 , \6675 , \6687 );
mnot \mul_7_15_g34651/U$4 ( \6689 , \6688 );
mor \mul_7_15_g34651/U$2 ( \6690 , \6658 , \6689 );
mnot \mul_7_15_g35279/U$3 ( \6691 , \6492 );
mnot \mul_7_15_g35730/U$3 ( \6692 , \4066 );
mnot \mul_7_15_g35730/U$4 ( \6693 , \6541 );
mor \mul_7_15_g35730/U$2 ( \6694 , \6692 , \6693 );
mnand \mul_7_15_g35804/U$1 ( \6695 , \5433 , \4519 );
mnand \mul_7_15_g35730/U$1 ( \6696 , \6694 , \6695 );
mnot \mul_7_15_g35279/U$4 ( \6697 , \6696 );
mor \mul_7_15_g35279/U$2 ( \6698 , \6691 , \6697 );
mnand \mul_7_15_g35442/U$1 ( \6699 , \6665 , \5266 );
mnand \mul_7_15_g35279/U$1 ( \6700 , \6698 , \6699 );
mnot \mul_7_15_g34780/U$3 ( \6701 , \6700 );
mand \mul_7_15_g35673/U$2 ( \6702 , \4079 , \4917 );
mnot \mul_7_15_g35673/U$4 ( \6703 , \4079 );
mand \mul_7_15_g35673/U$3 ( \6704 , \6703 , \4732 );
mnor \mul_7_15_g35673/U$1 ( \6705 , \6702 , \6704 );
mnot \mul_7_15_g35155/U$3 ( \6706 , \6705 );
mnot \mul_7_15_g35155/U$4 ( \6707 , \4632 );
mor \mul_7_15_g35155/U$2 ( \6708 , \6706 , \6707 );
mnot \mul_7_15_g35722/U$3 ( \6709 , \4076 );
mnot \mul_7_15_g35722/U$4 ( \6710 , \4535 );
mor \mul_7_15_g35722/U$2 ( \6711 , \6709 , \6710 );
mnand \mul_7_15_g37185/U$1 ( \6712 , \4917 , \5284 );
mnand \mul_7_15_g35722/U$1 ( \6713 , \6711 , \6712 );
mnand \mul_7_15_g35464/U$1 ( \6714 , \4453 , \6713 );
mnand \mul_7_15_g35155/U$1 ( \6715 , \6708 , \6714 );
mnot \mul_7_15_g34780/U$4 ( \6716 , \6715 );
mor \mul_7_15_g34780/U$2 ( \6717 , \6701 , \6716 );
mnot \mul_7_15_g35154/U$1 ( \6718 , \6715 );
mnot \g37275/U$3 ( \6719 , \6718 );
mnot \mul_7_15_g35278/U$1 ( \6720 , \6700 );
mnot \g37275/U$4 ( \6721 , \6720 );
mor \g37275/U$2 ( \6722 , \6719 , \6721 );
mnot \mul_7_15_g35745/U$3 ( \6723 , \4098 );
mnot \mul_7_15_g35745/U$4 ( \6724 , \4493 );
mor \mul_7_15_g35745/U$2 ( \6725 , \6723 , \6724 );
mnand \mul_7_15_g35900/U$1 ( \6726 , \4285 , \5418 );
mnand \mul_7_15_g35745/U$1 ( \6727 , \6725 , \6726 );
mnot \mul_7_15_g35111/U$3 ( \6728 , \6727 );
mnot \mul_7_15_g35111/U$4 ( \6729 , \4430 );
mor \mul_7_15_g35111/U$2 ( \6730 , \6728 , \6729 );
mnot \mul_7_15_g35664/U$3 ( \6731 , \4082 );
mnot \mul_7_15_g35664/U$4 ( \6732 , \4493 );
mor \mul_7_15_g35664/U$2 ( \6733 , \6731 , \6732 );
mnand \mul_7_15_g35886/U$1 ( \6734 , \4283 , \5526 );
mnand \mul_7_15_g35664/U$1 ( \6735 , \6733 , \6734 );
mnand \mul_7_15_g35369/U$1 ( \6736 , \6735 , \5160 );
mnand \mul_7_15_g35111/U$1 ( \6737 , \6730 , \6736 );
mnand \g37275/U$1 ( \6738 , \6722 , \6737 );
mnand \mul_7_15_g34780/U$1 ( \6739 , \6717 , \6738 );
mnand \mul_7_15_g34651/U$1 ( \6740 , \6690 , \6739 );
mnot \mul_7_15_g34819/U$1 ( \6741 , \6688 );
mnot \mul_7_15_g34927/U$1 ( \6742 , \6657 );
mnand \mul_7_15_g34735/U$1 ( \6743 , \6741 , \6742 );
mnand \mul_7_15_g34624/U$1 ( \6744 , \6740 , \6743 );
mnot \mul_7_15_g34605/U$1 ( \6745 , \6744 );
mnot \mul_7_15_g34550/U$4 ( \6746 , \6745 );
mor \mul_7_15_g34550/U$2 ( \6747 , \6635 , \6746 );
mnot \mul_7_15_g34555/U$2 ( \6748 , \6634 );
mnand \mul_7_15_g34555/U$1 ( \6749 , \6748 , \6744 );
mnand \mul_7_15_g34550/U$1 ( \6750 , \6747 , \6749 );
mnand \mul_7_15_g35011/U$1 ( \6751 , \6673 , \6659 );
mnot \mul_7_15_g34883/U$3 ( \6752 , \6751 );
mnot \mul_7_15_g34883/U$4 ( \6753 , \6686 );
mor \mul_7_15_g34883/U$2 ( \6754 , \6752 , \6753 );
mnand \mul_7_15_g35012/U$1 ( \6755 , \6670 , \6660 );
mnand \mul_7_15_g34883/U$1 ( \6756 , \6754 , \6755 );
mnot \mul_7_15_g35698/U$3 ( \6757 , \4026 );
mnot \mul_7_15_g35698/U$4 ( \6758 , \5301 );
mor \mul_7_15_g35698/U$2 ( \6759 , \6757 , \6758 );
mnand \mul_7_15_g35845/U$1 ( \6760 , \4616 , \4969 );
mnand \mul_7_15_g35698/U$1 ( \6761 , \6759 , \6760 );
mnot \mul_7_15_g35100/U$3 ( \6762 , \6761 );
mnot \mul_7_15_g35100/U$4 ( \6763 , \4611 );
mor \mul_7_15_g35100/U$2 ( \6764 , \6762 , \6763 );
mnot \mul_7_15_g35720/U$3 ( \6765 , \4021 );
mnot \mul_7_15_g35720/U$4 ( \6766 , \5138 );
mor \mul_7_15_g35720/U$2 ( \6767 , \6765 , \6766 );
mnand \mul_7_15_g35872/U$1 ( \6768 , \4745 , \4780 );
mnand \mul_7_15_g35720/U$1 ( \6769 , \6767 , \6768 );
mnand \mul_7_15_g35341/U$1 ( \6770 , \4881 , \6769 );
mnand \mul_7_15_g35100/U$1 ( \6771 , \6764 , \6770 );
mnot \mul_7_15_g35099/U$1 ( \6772 , \6771 );
mnot \mul_7_15_g34938/U$3 ( \6773 , \6772 );
mand \mul_7_15_g35097/U$2 ( \6774 , \4632 , \6713 );
mand \mul_7_15_g35097/U$3 ( \6775 , \4453 , \6607 );
mnor \mul_7_15_g35097/U$1 ( \6776 , \6774 , \6775 );
mnot \mul_7_15_g34938/U$4 ( \6777 , \6776 );
mor \mul_7_15_g34938/U$2 ( \6778 , \6773 , \6777 );
mnot \mul_7_15_g35098/U$3 ( \6779 , \6735 );
mnot \mul_7_15_g35098/U$4 ( \6780 , \4338 );
mor \mul_7_15_g35098/U$2 ( \6781 , \6779 , \6780 );
mnand \mul_7_15_g35386/U$1 ( \6782 , \6628 , \4341 );
mnand \mul_7_15_g35098/U$1 ( \6783 , \6781 , \6782 );
mnand \mul_7_15_g34938/U$1 ( \6784 , \6778 , \6783 );
mnot \mul_7_15_g36403/U$2 ( \6785 , \6776 );
mnand \mul_7_15_g36403/U$1 ( \6786 , \6785 , \6771 );
mnand \mul_7_15_g34909/U$1 ( \6787 , \6784 , \6786 );
mxor \mul_7_15_g34542/U$1 ( \6788 , \6756 , \6787 );
mnot \mul_7_15_g35108/U$3 ( \6789 , \6769 );
mnot \mul_7_15_g35108/U$4 ( \6790 , \4610 );
mor \mul_7_15_g35108/U$2 ( \6791 , \6789 , \6790 );
mnot \mul_7_15_g35651/U$3 ( \6792 , \4017 );
mnot \mul_7_15_g35651/U$4 ( \6793 , \5138 );
mor \mul_7_15_g35651/U$2 ( \6794 , \6792 , \6793 );
mnand \mul_7_15_g35842/U$1 ( \6795 , \4745 , \4662 );
mnand \mul_7_15_g35651/U$1 ( \6796 , \6794 , \6795 );
mnand \mul_7_15_g35354/U$1 ( \6797 , \6796 , \5146 );
mnand \mul_7_15_g35108/U$1 ( \6798 , \6791 , \6797 );
mnor \mul_7_15_g35752/U$1 ( \6799 , \4098 , \3573 );
mnot \mul_7_15_g35498/U$3 ( \6800 , \6799 );
mnot \mul_7_15_g35498/U$4 ( \6801 , \4284 );
mand \mul_7_15_g35498/U$2 ( \6802 , \6800 , \6801 );
mnot \mul_7_15_g35528/U$3 ( \6803 , \4098 );
mnot \mul_7_15_g35528/U$4 ( \6804 , \3573 );
mor \mul_7_15_g35528/U$2 ( \6805 , \6803 , \6804 );
mnand \mul_7_15_g35528/U$1 ( \6806 , \6805 , \4154 );
mnor \mul_7_15_g35498/U$1 ( \6807 , \6802 , \6806 );
mnot \mul_7_15_g34957/U$3 ( \6808 , \6807 );
mor \mul_7_15_g35021/U$2 ( \6809 , \6180 , \4862 );
mnand \mul_7_15_g35266/U$1 ( \6810 , \4862 , \6684 , \4858 );
mnand \mul_7_15_g35021/U$1 ( \6811 , \6809 , \6810 );
mnot \mul_7_15_g35020/U$1 ( \6812 , \6811 );
mnot \mul_7_15_g34957/U$4 ( \6813 , \6812 );
mor \mul_7_15_g34957/U$2 ( \6814 , \6808 , \6813 );
mor \mul_7_15_g34957/U$5 ( \6815 , \6812 , \6807 );
mnand \mul_7_15_g34957/U$1 ( \6816 , \6814 , \6815 );
mxor \mul_7_15_g34660/U$1 ( \6817 , \6798 , \6816 );
mnot \mul_7_15_g35746/U$3 ( \6818 , \4098 );
mnot \mul_7_15_g35746/U$4 ( \6819 , \4163 );
mor \mul_7_15_g35746/U$2 ( \6820 , \6818 , \6819 );
mnand \mul_7_15_g35903/U$1 ( \6821 , \4170 , \5418 );
mnand \mul_7_15_g35746/U$1 ( \6822 , \6820 , \6821 );
mnot \mul_7_15_g35089/U$3 ( \6823 , \6822 );
mnot \mul_7_15_g35089/U$4 ( \6824 , \4159 );
mor \mul_7_15_g35089/U$2 ( \6825 , \6823 , \6824 );
mnand \mul_7_15_g35358/U$1 ( \6826 , \4317 , \6211 );
mnand \mul_7_15_g35089/U$1 ( \6827 , \6825 , \6826 );
mxor \mul_7_15_g34660/U$1_r1 ( \6828 , \6817 , \6827 );
mxor \mul_7_15_g34542/U$1_r1 ( \6829 , \6788 , \6828 );
mnot \mul_7_15_g34540/U$1 ( \6830 , \6829 );
mand \mul_7_15_g34483/U$2 ( \6831 , \6750 , \6830 );
mnot \mul_7_15_g34483/U$4 ( \6832 , \6750 );
mand \mul_7_15_g34483/U$3 ( \6833 , \6832 , \6829 );
mnor \mul_7_15_g34483/U$1 ( \6834 , \6831 , \6833 );
mnot \mul_7_15_g35696/U$3 ( \6835 , \4072 );
mnot \mul_7_15_g35696/U$4 ( \6836 , \5138 );
mor \mul_7_15_g35696/U$2 ( \6837 , \6835 , \6836 );
mnand \mul_7_15_g35822/U$1 ( \6838 , \4616 , \5089 );
mnand \mul_7_15_g35696/U$1 ( \6839 , \6837 , \6838 );
mnot \mul_7_15_g35085/U$3 ( \6840 , \6839 );
mnot \mul_7_15_g35085/U$4 ( \6841 , \4611 );
mor \mul_7_15_g35085/U$2 ( \6842 , \6840 , \6841 );
mnand \mul_7_15_g35356/U$1 ( \6843 , \4754 , \6761 );
mnand \mul_7_15_g35085/U$1 ( \6844 , \6842 , \6843 );
mbuf \mul_7_15_g35084/U$1 ( \6845 , \6844 );
mnot \mul_7_15_g34684/U$3 ( \6846 , \6845 );
mnot \mul_7_15_g34959/U$3 ( \6847 , \6656 );
mnot \mul_7_15_g35023/U$1 ( \6848 , \6650 );
mnot \mul_7_15_g34959/U$4 ( \6849 , \6848 );
mor \mul_7_15_g34959/U$2 ( \6850 , \6847 , \6849 );
mnot \mul_7_15_g34977/U$2 ( \6851 , \6656 );
mnand \mul_7_15_g34977/U$1 ( \6852 , \6851 , \6650 );
mnand \mul_7_15_g34959/U$1 ( \6853 , \6850 , \6852 );
mbuf \mul_7_15_g34926/U$1 ( \6854 , \6853 );
mnot \mul_7_15_g34684/U$4 ( \6855 , \6854 );
mor \mul_7_15_g34684/U$2 ( \6856 , \6846 , \6855 );
mor \mul_7_15_g34718/U$2 ( \6857 , \6854 , \6845 );
mnand \mul_7_15_g35479/U$1 ( \6858 , \4800 , \4098 );
mnot \mul_7_15_g35478/U$1 ( \6859 , \6858 );
mnot \mul_7_15_g34777/U$3 ( \6860 , \6859 );
mnand \mul_7_15_g35305/U$1 ( \6861 , \6382 , \4859 );
mor \mul_7_15_g35017/U$2 ( \6862 , \6861 , \4948 );
mnand \mul_7_15_g35381/U$1 ( \6863 , \4863 , \6646 );
mnand \mul_7_15_g35017/U$1 ( \6864 , \6862 , \6863 );
mnot \mul_7_15_g34777/U$4 ( \6865 , \6864 );
mor \mul_7_15_g34777/U$2 ( \6866 , \6860 , \6865 );
mor \mul_7_15_g34874/U$2 ( \6867 , \6864 , \6859 );
mnot \mul_7_15_g35195/U$3 ( \6868 , \6423 );
mnot \mul_7_15_g35195/U$4 ( \6869 , \4632 );
mor \mul_7_15_g35195/U$2 ( \6870 , \6868 , \6869 );
mnand \mul_7_15_g35418/U$1 ( \6871 , \4453 , \6705 );
mnand \mul_7_15_g35195/U$1 ( \6872 , \6870 , \6871 );
mnand \mul_7_15_g34874/U$1 ( \6873 , \6867 , \6872 );
mnand \mul_7_15_g34777/U$1 ( \6874 , \6866 , \6873 );
mnand \mul_7_15_g34718/U$1 ( \6875 , \6857 , \6874 );
mnand \mul_7_15_g34684/U$1 ( \6876 , \6856 , \6875 );
mnot \mul_7_15_g34672/U$1 ( \6877 , \6876 );
mnot \mul_7_15_g34965/U$3 ( \6878 , \6783 );
mnot \mul_7_15_g34965/U$4 ( \6879 , \6772 );
mor \mul_7_15_g34965/U$2 ( \6880 , \6878 , \6879 );
mor \mul_7_15_g34965/U$5 ( \6881 , \6783 , \6772 );
mnand \mul_7_15_g34965/U$1 ( \6882 , \6880 , \6881 );
mbuf \mul_7_15_g35096/U$1 ( \6883 , \6776 );
mnot \mul_7_15_g35095/U$1 ( \6884 , \6883 );
mand \mul_7_15_g34892/U$2 ( \6885 , \6882 , \6884 );
mnot \mul_7_15_g34892/U$4 ( \6886 , \6882 );
mand \mul_7_15_g34892/U$3 ( \6887 , \6886 , \6883 );
mnor \mul_7_15_g34892/U$1 ( \6888 , \6885 , \6887 );
mnot \mul_7_15_g34850/U$1 ( \6889 , \6888 );
mnand \mul_7_15_g34611/U$1 ( \6890 , \6877 , \6889 );
mnot \mul_7_15_g34511/U$3 ( \6891 , \6890 );
mnot \mul_7_15_g34725/U$3 ( \6892 , \6742 );
mnot \mul_7_15_g34725/U$4 ( \6893 , \6688 );
mor \mul_7_15_g34725/U$2 ( \6894 , \6892 , \6893 );
mnand \mul_7_15_g34734/U$1 ( \6895 , \6741 , \6657 );
mnand \mul_7_15_g34725/U$1 ( \6896 , \6894 , \6895 );
mand \mul_7_15_g34632/U$2 ( \6897 , \6896 , \6739 );
mnot \mul_7_15_g34632/U$4 ( \6898 , \6896 );
mnot \mul_7_15_g34776/U$1 ( \6899 , \6739 );
mand \mul_7_15_g34632/U$3 ( \6900 , \6898 , \6899 );
mnor \mul_7_15_g34632/U$1 ( \6901 , \6897 , \6900 );
mnot \mul_7_15_g34511/U$4 ( \6902 , \6901 );
mor \mul_7_15_g34511/U$2 ( \6903 , \6891 , \6902 );
mnot \mul_7_15_g36377/U$2 ( \6904 , \6877 );
mnand \mul_7_15_g36377/U$1 ( \6905 , \6904 , \6888 );
mnand \mul_7_15_g34511/U$1 ( \6906 , \6903 , \6905 );
mnot \mul_7_15_g34500/U$1 ( \6907 , \6906 );
mnand \mul_7_15_g34421/U$1 ( \6908 , \6834 , \6907 );
mxor \mul_7_15_g34852/U$1 ( \6909 , \6700 , \6737 );
mxnor \mul_7_15_g34852/U$1_r1 ( \6910 , \6909 , \6715 );
mnand \mul_7_15_g35003/U$1 ( \6911 , \6384 , \6372 );
mnot \mul_7_15_g34879/U$2 ( \6912 , \6911 );
mnot \mul_7_15_g35149/U$3 ( \6913 , \6410 );
mnot \mul_7_15_g35149/U$4 ( \6914 , \4611 );
mor \mul_7_15_g35149/U$2 ( \6915 , \6913 , \6914 );
mnand \mul_7_15_g35460/U$1 ( \6916 , \6839 , \4754 );
mnand \mul_7_15_g35149/U$1 ( \6917 , \6915 , \6916 );
mnot \mul_7_15_g35298/U$3 ( \6918 , \6401 );
mnot \mul_7_15_g35298/U$4 ( \6919 , \6492 );
mor \mul_7_15_g35298/U$2 ( \6920 , \6918 , \6919 );
mnand \mul_7_15_g35431/U$1 ( \6921 , \6696 , \5266 );
mnand \mul_7_15_g35298/U$1 ( \6922 , \6920 , \6921 );
mor \mul_7_15_g36409/U$1 ( \6923 , \6917 , \6922 );
mnand \mul_7_15_g34879/U$1 ( \6924 , \6912 , \6923 );
mnand \mul_7_15_g34996/U$1 ( \6925 , \6917 , \6922 );
mand \mul_7_15_g34783/U$1 ( \6926 , \6924 , \6925 );
mxor \mul_7_15_g34548/U$1 ( \6927 , \6910 , \6926 );
mxor \mul_7_15_g34702/U$1 ( \6928 , \6844 , \6853 );
mxnor \mul_7_15_g34702/U$1_r1 ( \6929 , \6928 , \6874 );
mxor \mul_7_15_g34548/U$1_r1 ( \6930 , \6927 , \6929 );
mxor \mul_7_15_g34793/U$1 ( \6931 , \6858 , \6864 );
mxnor \mul_7_15_g34793/U$1_r1 ( \6932 , \6931 , \6872 );
mxor \mul_7_15_g34812/U$4 ( \6933 , \6403 , \6412 );
mand \mul_7_15_g34812/U$3 ( \6934 , \6933 , \6426 );
mand \mul_7_15_g34812/U$5 ( \6935 , \6403 , \6412 );
mor \mul_7_15_g34812/U$2 ( \6936 , \6934 , \6935 );
mxor \mul_7_15_g34602/U$4 ( \6937 , \6932 , \6936 );
mxor \mul_7_15_g34796/U$1 ( \6938 , \6922 , \6917 );
mxnor \mul_7_15_g34796/U$1_r1 ( \6939 , \6938 , \6911 );
mand \mul_7_15_g34602/U$3 ( \6940 , \6937 , \6939 );
mand \mul_7_15_g34602/U$5 ( \6941 , \6932 , \6936 );
mor \mul_7_15_g34602/U$2 ( \6942 , \6940 , \6941 );
mnot \mul_7_15_g34601/U$1 ( \6943 , \6942 );
mnand \mul_7_15_g34505/U$1 ( \6944 , \6930 , \6943 );
mxor \mul_7_15_g34602/U$1 ( \6945 , \6932 , \6936 );
mxor \mul_7_15_g34602/U$1_r1 ( \6946 , \6945 , \6939 );
mnot \mul_7_15_g34600/U$1 ( \6947 , \6946 );
mxor \mul_7_15_g34594/U$4 ( \6948 , \6388 , \6392 );
mand \mul_7_15_g34594/U$3 ( \6949 , \6948 , \6427 );
mand \mul_7_15_g34594/U$5 ( \6950 , \6388 , \6392 );
mor \mul_7_15_g34594/U$2 ( \6951 , \6949 , \6950 );
mnot \mul_7_15_g34593/U$1 ( \6952 , \6951 );
mnand \mul_7_15_g34560/U$1 ( \6953 , \6947 , \6952 );
mand \mul_7_15_g34488/U$1 ( \6954 , \6944 , \6953 );
mand \mul_7_15_g34606/U$2 ( \6955 , \6876 , \6888 );
mnot \mul_7_15_g34606/U$4 ( \6956 , \6876 );
mand \mul_7_15_g34606/U$3 ( \6957 , \6956 , \6889 );
mnor \mul_7_15_g34606/U$1 ( \6958 , \6955 , \6957 );
mxnor \mul_7_15_g36372/U$1 ( \6959 , \6958 , \6901 );
mxor \mul_7_15_g34548/U$4 ( \6960 , \6910 , \6926 );
mand \mul_7_15_g34548/U$3 ( \6961 , \6960 , \6929 );
mand \mul_7_15_g34548/U$5 ( \6962 , \6910 , \6926 );
mor \mul_7_15_g34548/U$2 ( \6963 , \6961 , \6962 );
mnand \mul_7_15_g34459/U$1 ( \6964 , \6959 , \6963 );
mnand \mul_7_15_g34384/U$1 ( \6965 , \6908 , \6954 , \6964 );
mnot \mul_7_15_g34383/U$1 ( \6966 , \6965 );
mnot \mul_7_15_g34344/U$4 ( \6967 , \6966 );
mor \mul_7_15_g34344/U$2 ( \6968 , \6602 , \6967 );
mnot \g37055/U$2 ( \6969 , \6834 );
mnand \g37055/U$1 ( \6970 , \6969 , \6906 );
mnot \mul_7_15_g34499/U$1 ( \6971 , \6959 );
mnot \mul_7_15_g34547/U$1 ( \6972 , \6963 );
mnand \mul_7_15_g34461/U$1 ( \6973 , \6971 , \6972 );
mnand \mul_7_15_g34397/U$1 ( \6974 , \6970 , \6973 );
mnot \mul_7_15_g34546/U$1 ( \6975 , \6930 );
mnand \mul_7_15_g34508/U$1 ( \6976 , \6975 , \6942 );
mnand \mul_7_15_g34556/U$1 ( \6977 , \6946 , \6951 );
mnand \mul_7_15_g34487/U$1 ( \6978 , \6976 , \6977 );
mand \mul_7_15_g34429/U$1 ( \6979 , \6964 , \6978 , \6944 );
mor \mul_7_15_g34366/U$2 ( \6980 , \6974 , \6979 );
mbuf \mul_7_15_g34420/U$1 ( \6981 , \6908 );
mnand \mul_7_15_g34366/U$1 ( \6982 , \6980 , \6981 );
mnand \mul_7_15_g34344/U$1 ( \6983 , \6968 , \6982 );
mxor \mul_7_15_g34854/U$1 ( \6984 , \6062 , \6088 );
mxnor \mul_7_15_g34854/U$1_r1 ( \6985 , \6984 , \6074 );
mnot \mul_7_15_g34779/U$3 ( \6986 , \6622 );
mnot \mul_7_15_g34779/U$4 ( \6987 , \6612 );
mor \mul_7_15_g34779/U$2 ( \6988 , \6986 , \6987 );
mor \mul_7_15_g34871/U$2 ( \6989 , \6612 , \6622 );
mnand \mul_7_15_g34871/U$1 ( \6990 , \6989 , \6633 );
mnand \mul_7_15_g34779/U$1 ( \6991 , \6988 , \6990 );
mnot \mul_7_15_g35128/U$3 ( \6992 , \6796 );
mnot \mul_7_15_g35128/U$4 ( \6993 , \4611 );
mor \mul_7_15_g35128/U$2 ( \6994 , \6992 , \6993 );
mnand \mul_7_15_g35419/U$1 ( \6995 , \4754 , \6108 );
mnand \mul_7_15_g35128/U$1 ( \6996 , \6994 , \6995 );
mnot \mul_7_15_g35127/U$1 ( \6997 , \6996 );
mnot \mul_7_15_g36398/U$2 ( \6998 , \6812 );
mnand \mul_7_15_g36398/U$1 ( \6999 , \6998 , \6807 );
mnand \mul_7_15_g34863/U$1 ( \7000 , \6997 , \6999 );
mand \mul_7_15_g34681/U$2 ( \7001 , \6991 , \7000 );
mnor \mul_7_15_g34862/U$1 ( \7002 , \6997 , \6999 );
mnor \mul_7_15_g34681/U$1 ( \7003 , \7001 , \7002 );
mxor \mul_7_15_g34567/U$1 ( \7004 , \6985 , \7003 );
mnot \mul_7_15_g35141/U$1 ( \7005 , \6113 );
mxor \g37154/U$1 ( \7006 , \6124 , \7005 );
mand \g37153/U$2 ( \7007 , \7006 , \6103 );
mnot \g37153/U$4 ( \7008 , \7006 );
mnot \mul_7_15_g35136/U$1 ( \7009 , \6103 );
mand \g37153/U$3 ( \7010 , \7008 , \7009 );
mnor \g37153/U$1 ( \7011 , \7007 , \7010 );
mxor \mul_7_15_g34567/U$1_r1 ( \7012 , \7004 , \7011 );
mnot \mul_7_15_g34566/U$1 ( \7013 , \7012 );
mnot \g37142/U$3 ( \7014 , \7013 );
mxor \g36481/U$1 ( \7015 , \6162 , \6192 );
mxnor \g36481/U$1_r1 ( \7016 , \7015 , \6232 );
mnot \g37142/U$4 ( \7017 , \7016 );
mor \g37142/U$2 ( \7018 , \7014 , \7017 );
mnot \mul_7_15_g34585/U$1 ( \7019 , \7016 );
mnot \g37143/U$3 ( \7020 , \7019 );
mnot \g37143/U$4 ( \7021 , \7012 );
mor \g37143/U$2 ( \7022 , \7020 , \7021 );
mxor \mul_7_15_g34886/U$1 ( \7023 , \6173 , \6175 );
mxor \mul_7_15_g34886/U$1_r1 ( \7024 , \7023 , \6186 );
mnot \mul_7_15_g34529/U$3 ( \7025 , \7024 );
mxor \mul_7_15_g34660/U$4 ( \7026 , \6798 , \6816 );
mand \mul_7_15_g34660/U$3 ( \7027 , \7026 , \6827 );
mand \mul_7_15_g34660/U$5 ( \7028 , \6798 , \6816 );
mor \mul_7_15_g34660/U$2 ( \7029 , \7027 , \7028 );
mnot \mul_7_15_g34659/U$1 ( \7030 , \7029 );
mnot \mul_7_15_g34529/U$4 ( \7031 , \7030 );
mor \mul_7_15_g34529/U$2 ( \7032 , \7025 , \7031 );
mnot \mul_7_15_g34968/U$3 ( \7033 , \6229 );
mnot \mul_7_15_g34968/U$4 ( \7034 , \6205 );
mor \mul_7_15_g34968/U$2 ( \7035 , \7033 , \7034 );
mor \mul_7_15_g34968/U$5 ( \7036 , \6205 , \6229 );
mnand \mul_7_15_g34968/U$1 ( \7037 , \7035 , \7036 );
mand \mul_7_15_g34894/U$2 ( \7038 , \7037 , \6216 );
mnot \mul_7_15_g34894/U$4 ( \7039 , \7037 );
mand \mul_7_15_g34894/U$3 ( \7040 , \7039 , \6217 );
mnor \mul_7_15_g34894/U$1 ( \7041 , \7038 , \7040 );
mnand \mul_7_15_g34529/U$1 ( \7042 , \7032 , \7041 );
mnot \mul_7_15_g36394/U$2 ( \7043 , \7024 );
mnand \mul_7_15_g36394/U$1 ( \7044 , \7043 , \7029 );
mnand \mul_7_15_g34512/U$1 ( \7045 , \7042 , \7044 );
mnand \g37143/U$1 ( \7046 , \7022 , \7045 );
mnand \g37142/U$1 ( \7047 , \7018 , \7046 );
mnot \mul_7_15_g36360/U$2 ( \7048 , \7047 );
mxor \g36485/U$1 ( \7049 , \6090 , \6051 );
mnot \mul_7_15_g34809/U$1 ( \7050 , \6127 );
mand \mul_7_15_g34609/U$2 ( \7051 , \7049 , \7050 );
mnot \mul_7_15_g34609/U$4 ( \7052 , \7049 );
mand \mul_7_15_g34609/U$3 ( \7053 , \7052 , \6127 );
mnor \mul_7_15_g34609/U$1 ( \7054 , \7051 , \7053 );
mxor \mul_7_15_g34567/U$4 ( \7055 , \6985 , \7003 );
mand \mul_7_15_g34567/U$3 ( \7056 , \7055 , \7011 );
mand \mul_7_15_g34567/U$5 ( \7057 , \6985 , \7003 );
mor \mul_7_15_g34567/U$2 ( \7058 , \7056 , \7057 );
mxor \mul_7_15_g34414/U$1 ( \7059 , \7054 , \7058 );
mand \mul_7_15_g34607/U$2 ( \7060 , \6251 , \6261 );
mnot \mul_7_15_g34607/U$4 ( \7061 , \6251 );
mnot \mul_7_15_g34664/U$1 ( \7062 , \6261 );
mand \mul_7_15_g34607/U$3 ( \7063 , \7061 , \7062 );
mnor \mul_7_15_g34607/U$1 ( \7064 , \7060 , \7063 );
mxor \g36785/U$1 ( \7065 , \6236 , \7064 );
mxor \mul_7_15_g34414/U$1_r1 ( \7066 , \7059 , \7065 );
mbuf \mul_7_15_g34412/U$1 ( \7067 , \7066 );
mnand \mul_7_15_g36360/U$1 ( \7068 , \7048 , \7067 );
mxor \mul_7_15_g34374/U$1 ( \7069 , \6161 , \6267 );
mxor \mul_7_15_g34374/U$1_r1 ( \7070 , \7069 , \6270 );
mnot \mul_7_15_g34339/U$2 ( \7071 , \7070 );
mxor \mul_7_15_g34414/U$4 ( \7072 , \7054 , \7058 );
mand \mul_7_15_g34414/U$3 ( \7073 , \7072 , \7065 );
mand \mul_7_15_g34414/U$5 ( \7074 , \7054 , \7058 );
mor \mul_7_15_g34414/U$2 ( \7075 , \7073 , \7074 );
mnand \mul_7_15_g34339/U$1 ( \7076 , \7071 , \7075 );
mxor \mul_7_15_g2/U$1 ( \7077 , \7016 , \7045 );
mand \mul_7_15_g34415/U$2 ( \7078 , \7077 , \7012 );
mnot \mul_7_15_g34415/U$4 ( \7079 , \7077 );
mand \mul_7_15_g34415/U$3 ( \7080 , \7079 , \7013 );
mnor \mul_7_15_g34415/U$1 ( \7081 , \7078 , \7080 );
mnot \mul_7_15_g34921/U$1 ( \7082 , \6999 );
mnot \mul_7_15_g34789/U$3 ( \7083 , \7082 );
mnot \mul_7_15_g34789/U$4 ( \7084 , \6997 );
mor \mul_7_15_g34789/U$2 ( \7085 , \7083 , \7084 );
mor \mul_7_15_g34789/U$5 ( \7086 , \6997 , \7082 );
mnand \mul_7_15_g34789/U$1 ( \7087 , \7085 , \7086 );
mxor \g36764/U$1 ( \7088 , \6991 , \7087 );
mbuf \mul_7_15_g34661/U$1 ( \7089 , \7088 );
mnot \mul_7_15_g34465/U$2 ( \7090 , \7089 );
mxor \mul_7_15_g34519/U$1 ( \7091 , \7024 , \7029 );
mxnor \mul_7_15_g34519/U$1_r1 ( \7092 , \7091 , \7041 );
mnot \mul_7_15_g34494/U$1 ( \7093 , \7092 );
mnand \mul_7_15_g34465/U$1 ( \7094 , \7090 , \7093 );
mxor \mul_7_15_g34542/U$4 ( \7095 , \6756 , \6787 );
mand \mul_7_15_g34542/U$3 ( \7096 , \7095 , \6828 );
mand \mul_7_15_g34542/U$5 ( \7097 , \6756 , \6787 );
mor \mul_7_15_g34542/U$2 ( \7098 , \7096 , \7097 );
mbuf \mul_7_15_g34541/U$1 ( \7099 , \7098 );
mand \mul_7_15_g34430/U$2 ( \7100 , \7094 , \7099 );
mand \g37244/U$1 ( \7101 , \7092 , \7089 );
mnor \mul_7_15_g34430/U$1 ( \7102 , \7100 , \7101 );
mnand \mul_7_15_g34355/U$1 ( \7103 , \7081 , \7102 );
mnot \mul_7_15_g34471/U$3 ( \7104 , \6829 );
mnot \mul_7_15_g36380/U$2 ( \7105 , \6634 );
mnand \mul_7_15_g36380/U$1 ( \7106 , \7105 , \6745 );
mnot \mul_7_15_g34471/U$4 ( \7107 , \7106 );
mor \mul_7_15_g34471/U$2 ( \7108 , \7104 , \7107 );
mnand \mul_7_15_g34561/U$1 ( \7109 , \6744 , \6634 );
mnand \mul_7_15_g34471/U$1 ( \7110 , \7108 , \7109 );
mnot \mul_7_15_g36368/U$2 ( \7111 , \7110 );
mxor \mul_7_15_g34456/U$1 ( \7112 , \7088 , \7098 );
mxnor \mul_7_15_g34456/U$1_r1 ( \7113 , \7112 , \7092 );
mnand \mul_7_15_g36368/U$1 ( \7114 , \7111 , \7113 );
mand \mul_7_15_g36347/U$1 ( \7115 , \7103 , \7114 );
mand \mul_7_15_g34288/U$1 ( \7116 , \7068 , \7076 , \7115 );
mnand \mul_7_15_g34275/U$1 ( \7117 , \6983 , \7116 );
mnot \mul_7_15_g36365/U$2 ( \7118 , \7075 );
mnand \mul_7_15_g36365/U$1 ( \7119 , \7118 , \7070 );
mnot \mul_7_15_g34250/U$3 ( \7120 , \7119 );
mnot \mul_7_15_g34341/U$2 ( \7121 , \7103 );
mnot \mul_7_15_g36364/U$2 ( \7122 , \7113 );
mnand \mul_7_15_g36364/U$1 ( \7123 , \7122 , \7110 );
mnor \mul_7_15_g34341/U$1 ( \7124 , \7121 , \7123 );
mnot \mul_7_15_g34386/U$1 ( \7125 , \7081 );
mnot \mul_7_15_g34411/U$1 ( \7126 , \7102 );
mnand \mul_7_15_g34359/U$1 ( \7127 , \7125 , \7126 );
mnot \mul_7_15_g34362/U$2 ( \7128 , \7066 );
mnand \mul_7_15_g34362/U$1 ( \7129 , \7128 , \7047 );
mnand \mul_7_15_g34343/U$1 ( \7130 , \7127 , \7129 );
mor \mul_7_15_g34285/U$2 ( \7131 , \7124 , \7130 );
mnand \mul_7_15_g34285/U$1 ( \7132 , \7131 , \7068 );
mnot \mul_7_15_g34250/U$4 ( \7133 , \7132 );
mor \mul_7_15_g34250/U$2 ( \7134 , \7120 , \7133 );
mbuf \mul_7_15_g34338/U$1 ( \7135 , \7076 );
mnand \mul_7_15_g34250/U$1 ( \7136 , \7134 , \7135 );
mnand \mul_7_15_g34232/U$1 ( \7137 , \7117 , \7136 );
mnand \mul_7_15_g34209/U$1 ( \7138 , \5707 , \6290 , \7137 );
mnot \mul_7_15_g34200/U$3 ( \7139 , \6288 );
mnand \mul_7_15_g34240/U$1 ( \7140 , \6044 , \6149 );
mnot \g36781/U$3 ( \7141 , \7140 );
mnand \mul_7_15_g34259/U$1 ( \7142 , \6276 , \6273 );
mnot \g36781/U$4 ( \7143 , \7142 );
mor \g36781/U$2 ( \7144 , \7141 , \7143 );
mnand \g36781/U$1 ( \7145 , \7144 , \6151 );
mor \mul_7_15_g34206/U$2 ( \7146 , \7145 , \6033 );
mnand \mul_7_15_g34241/U$1 ( \7147 , \5849 , \6032 );
mnand \mul_7_15_g34206/U$1 ( \7148 , \7146 , \7147 );
mnot \mul_7_15_g34200/U$4 ( \7149 , \7148 );
mor \mul_7_15_g34200/U$2 ( \7150 , \7139 , \7149 );
mnot \fopt36910/U$1 ( \7151 , \6287 );
mnot \mul_7_15_g34371/U$1 ( \7152 , \6281 );
mnand \mul_7_15_g34324/U$1 ( \7153 , \7151 , \7152 );
mnand \mul_7_15_g34200/U$1 ( \7154 , \7150 , \7153 );
mnand \mul_7_15_g34197/U$1 ( \7155 , \7154 , \5707 );
mbuf \mul_7_15_g34234/U$1 ( \7156 , \5649 );
mnot \mul_7_15_g34349/U$1 ( \7157 , \5651 );
mnot \mul_7_15_g34372/U$1 ( \7158 , \5705 );
mnand \mul_7_15_g34310/U$1 ( \7159 , \7157 , \7158 );
mor \mul_7_15_g36357/U$1 ( \7160 , \5354 , \5617 );
mnand \mul_7_15_g34260/U$1 ( \7161 , \7159 , \7160 );
mand \mul_7_15_g34213/U$2 ( \7162 , \7156 , \7161 );
mbuf \fopt36735/U$1 ( \7163 , \5648 );
mnot \fopt36734/U$1 ( \7164 , \7163 );
mor \mul_7_15_g36355/U$1 ( \7165 , \5640 , \5622 );
mor \mul_7_15_g34233/U$2 ( \7166 , \7164 , \7165 );
mor \mul_7_15_g36356/U$1 ( \7167 , \5647 , \5645 );
mnand \mul_7_15_g34233/U$1 ( \7168 , \7166 , \7167 );
mnor \mul_7_15_g34213/U$1 ( \7169 , \7162 , \7168 );
mnand \mul_7_15_g34194/U$1 ( \7170 , \7138 , \7155 , \7169 );
mnot \mul_7_15_g34187/U$4 ( \7171 , \7170 );
mor \mul_7_15_g34187/U$2 ( \7172 , \5071 , \7171 );
mnot \mul_7_15_g34521/U$1 ( \7173 , \5069 );
mnot \mul_7_15_g34202/U$3 ( \7174 , \7173 );
mnot \mul_7_15_g34208/U$3 ( \7175 , \5045 );
mnot \mul_7_15_g34222/U$3 ( \7176 , \4370 );
mnand \mul_7_15_g34330/U$1 ( \7177 , \4828 , \5003 );
mnor \mul_7_15_g34317/U$1 ( \7178 , \4825 , \7177 );
mand \mul_7_15_g34364/U$1 ( \7179 , \4822 , \4824 );
mnor \mul_7_15_g34292/U$1 ( \7180 , \7178 , \7179 );
mnand \mul_7_15_g34423/U$1 ( \7181 , \5010 , \5012 );
mnot \mul_7_15_g36366/U$2 ( \7182 , \7181 );
mand \mul_7_15_g34406/U$1 ( \7183 , \4488 , \4586 );
mnor \mul_7_15_g36366/U$1 ( \7184 , \7182 , \7183 );
mand \mul_7_15_g34252/U$2 ( \7185 , \7180 , \7184 );
mnot \g36780/U$3 ( \7186 , \4588 );
mnot \g36780/U$4 ( \7187 , \5013 );
mor \g36780/U$2 ( \7188 , \7186 , \7187 );
mnand \g36780/U$1 ( \7189 , \7188 , \7181 );
mnot \mul_7_15_g34334/U$1 ( \7190 , \7189 );
mnor \mul_7_15_g34252/U$1 ( \7191 , \7185 , \7190 );
mnot \mul_7_15_g34222/U$4 ( \7192 , \7191 );
mor \mul_7_15_g34222/U$2 ( \7193 , \7176 , \7192 );
mor \mul_7_15_g36369/U$1 ( \7194 , \4369 , \4293 );
mnand \mul_7_15_g34222/U$1 ( \7195 , \7193 , \7194 );
mnot \mul_7_15_g34208/U$4 ( \7196 , \7195 );
mor \mul_7_15_g34208/U$2 ( \7197 , \7175 , \7196 );
mnand \mul_7_15_g34462/U$1 ( \7198 , \5019 , \5044 );
mnand \mul_7_15_g34208/U$1 ( \7199 , \7197 , \7198 );
mnot \mul_7_15_g34202/U$4 ( \7200 , \7199 );
mor \mul_7_15_g34202/U$2 ( \7201 , \7174 , \7200 );
mnand \mul_7_15_g34525/U$1 ( \7202 , \5050 , \5068 );
mnand \mul_7_15_g34202/U$1 ( \7203 , \7201 , \7202 );
mnot \mul_7_15_g34201/U$1 ( \7204 , \7203 );
mnand \mul_7_15_g34187/U$1 ( \7205 , \7172 , \7204 );
mnot \mul_7_15_g35596/U$1 ( \7206 , \5064 );
mand \mul_7_15_g35247/U$2 ( \7207 , \4195 , \7206 );
mand \mul_7_15_g35247/U$3 ( \7208 , \4200 , \4253 );
mnor \mul_7_15_g35247/U$1 ( \7209 , \7207 , \7208 );
mnot \mul_7_15_g34949/U$3 ( \7210 , \7209 );
mnand \mul_7_15_g35774/U$1 ( \7211 , \4253 , \3997 );
mnot \mul_7_15_g34949/U$4 ( \7212 , \7211 );
mand \mul_7_15_g34949/U$2 ( \7213 , \7210 , \7212 );
mand \mul_7_15_g34949/U$5 ( \7214 , \7209 , \7211 );
mnor \mul_7_15_g34949/U$1 ( \7215 , \7213 , \7214 );
mnot \mul_7_15_g34726/U$3 ( \7216 , \7215 );
mxor \mul_7_15_g34832/U$4 ( \7217 , \5057 , \5059 );
mand \mul_7_15_g34832/U$3 ( \7218 , \7217 , \5066 );
mand \mul_7_15_g34832/U$5 ( \7219 , \5057 , \5059 );
mor \mul_7_15_g34832/U$2 ( \7220 , \7218 , \7219 );
mnot \mul_7_15_g34726/U$4 ( \7221 , \7220 );
mor \mul_7_15_g34726/U$2 ( \7222 , \7216 , \7221 );
mor \mul_7_15_g34726/U$5 ( \7223 , \7220 , \7215 );
mnand \mul_7_15_g34726/U$1 ( \7224 , \7222 , \7223 );
mnot \mul_7_15_g34538/U$3 ( \7225 , \7224 );
mxor \mul_7_15_g34599/U$4 ( \7226 , \5051 , \5055 );
mand \mul_7_15_g34599/U$3 ( \7227 , \7226 , \5067 );
mand \mul_7_15_g34599/U$5 ( \7228 , \5051 , \5055 );
mor \mul_7_15_g34599/U$2 ( \7229 , \7227 , \7228 );
mnot \mul_7_15_g34538/U$4 ( \7230 , \7229 );
mor \mul_7_15_g34538/U$2 ( \7231 , \7225 , \7230 );
mor \mul_7_15_g34538/U$5 ( \7232 , \7229 , \7224 );
mnand \mul_7_15_g34538/U$1 ( \7233 , \7231 , \7232 );
mnot \mul_7_15_g34537/U$1 ( \7234 , \7233 );
mand \mul_7_15_g34173/U$2 ( \7235 , \7205 , \7234 );
mnot \mul_7_15_g34173/U$4 ( \7236 , \7205 );
mand \mul_7_15_g34173/U$3 ( \7237 , \7236 , \7233 );
mnor \mul_7_15_g34173/U$1 ( \7238 , \7235 , \7237 );
mnot \fopt36702/U$1 ( \7239 , \5046 );
mnot \mul_7_15_g34185/U$3 ( \7240 , \7239 );
mnand \mul_7_15_g34195/U$1 ( \7241 , \7138 , \7155 , \7169 );
mnot \mul_7_15_g34185/U$4 ( \7242 , \7241 );
mor \mul_7_15_g34185/U$2 ( \7243 , \7240 , \7242 );
mnot \mul_7_15_g34207/U$1 ( \7244 , \7199 );
mnand \mul_7_15_g34185/U$1 ( \7245 , \7243 , \7244 );
mnand \mul_7_15_g34507/U$1 ( \7246 , \7173 , \7202 );
mnot \mul_7_15_g34506/U$1 ( \7247 , \7246 );
mand \mul_7_15_g34174/U$2 ( \7248 , \7245 , \7247 );
mnot \mul_7_15_g34174/U$4 ( \7249 , \7245 );
mand \mul_7_15_g34174/U$3 ( \7250 , \7249 , \7246 );
mnor \mul_7_15_g34174/U$1 ( \7251 , \7248 , \7250 );
mnot \mul_7_15_g34182/U$3 ( \7252 , \5015 );
mnot \mul_7_15_g34182/U$4 ( \7253 , \7241 );
mor \mul_7_15_g34182/U$2 ( \7254 , \7252 , \7253 );
mnot \mul_7_15_g34221/U$1 ( \7255 , \7195 );
mnand \mul_7_15_g34182/U$1 ( \7256 , \7254 , \7255 );
mnand \mul_7_15_g34442/U$1 ( \7257 , \5045 , \7198 );
mnot \mul_7_15_g34441/U$1 ( \7258 , \7257 );
mand \mul_7_15_g34175/U$2 ( \7259 , \7256 , \7258 );
mnot \mul_7_15_g34175/U$4 ( \7260 , \7256 );
mand \mul_7_15_g34175/U$3 ( \7261 , \7260 , \7257 );
mnor \mul_7_15_g34175/U$1 ( \7262 , \7259 , \7261 );
mnot \mul_7_15_g34266/U$1 ( \7263 , \5014 );
mnot \mul_7_15_g34186/U$3 ( \7264 , \7263 );
mnot \mul_7_15_g34186/U$4 ( \7265 , \7170 );
mor \mul_7_15_g34186/U$2 ( \7266 , \7264 , \7265 );
mnot \mul_7_15_g34251/U$1 ( \7267 , \7191 );
mnand \mul_7_15_g34186/U$1 ( \7268 , \7266 , \7267 );
mnand \mul_7_15_g34418/U$1 ( \7269 , \4370 , \7194 );
mnot \mul_7_15_g34417/U$1 ( \7270 , \7269 );
mand \mul_7_15_g34176/U$2 ( \7271 , \7268 , \7270 );
mnot \mul_7_15_g34176/U$4 ( \7272 , \7268 );
mand \mul_7_15_g34176/U$3 ( \7273 , \7272 , \7269 );
mnor \mul_7_15_g34176/U$1 ( \7274 , \7271 , \7273 );
mnot \mul_7_15_g34191/U$3 ( \7275 , \5006 );
mnot \mul_7_15_g34191/U$4 ( \7276 , \7170 );
mor \mul_7_15_g34191/U$2 ( \7277 , \7275 , \7276 );
mbuf \mul_7_15_g34291/U$1 ( \7278 , \7180 );
mnot \mul_7_15_g34290/U$1 ( \7279 , \7278 );
mand \mul_7_15_g34249/U$2 ( \7280 , \7279 , \4589 );
mnor \mul_7_15_g34249/U$1 ( \7281 , \7280 , \7183 );
mnand \mul_7_15_g34191/U$1 ( \7282 , \7277 , \7281 );
mnand \mul_7_15_g34396/U$1 ( \7283 , \5013 , \7181 );
mnot \mul_7_15_g34395/U$1 ( \7284 , \7283 );
mand \mul_7_15_g34177/U$2 ( \7285 , \7282 , \7284 );
mnot \mul_7_15_g34177/U$4 ( \7286 , \7282 );
mand \mul_7_15_g34177/U$3 ( \7287 , \7286 , \7283 );
mnor \mul_7_15_g34177/U$1 ( \7288 , \7285 , \7287 );
mnot \mul_7_15_g34318/U$1 ( \7289 , \5005 );
mnot \mul_7_15_g34181/U$3 ( \7290 , \7289 );
mnot \mul_7_15_g34181/U$4 ( \7291 , \7170 );
mor \mul_7_15_g34181/U$2 ( \7292 , \7290 , \7291 );
mnand \mul_7_15_g34181/U$1 ( \7293 , \7292 , \7278 );
mnot \mul_7_15_g36363/U$2 ( \7294 , \7183 );
mnand \mul_7_15_g36363/U$1 ( \7295 , \7294 , \4589 );
mnot \mul_7_15_g34377/U$1 ( \7296 , \7295 );
mand \mul_7_15_g34178/U$2 ( \7297 , \7293 , \7296 );
mnot \mul_7_15_g34178/U$4 ( \7298 , \7293 );
mand \mul_7_15_g34178/U$3 ( \7299 , \7298 , \7295 );
mnor \mul_7_15_g34178/U$1 ( \7300 , \7297 , \7299 );
mnot \mul_7_15_g34183/U$3 ( \7301 , \5004 );
mnot \mul_7_15_g34183/U$4 ( \7302 , \7241 );
mor \mul_7_15_g34183/U$2 ( \7303 , \7301 , \7302 );
mbuf \fopt36809/U$1 ( \7304 , \7177 );
mnand \mul_7_15_g34183/U$1 ( \7305 , \7303 , \7304 );
mor \mul_7_15_g36358/U$1 ( \7306 , \4825 , \7179 );
mnot \mul_7_15_g34325/U$1 ( \7307 , \7306 );
mand \mul_7_15_g34179/U$2 ( \7308 , \7305 , \7307 );
mnot \mul_7_15_g34179/U$4 ( \7309 , \7305 );
mand \mul_7_15_g34179/U$3 ( \7310 , \7309 , \7306 );
mnor \mul_7_15_g34179/U$1 ( \7311 , \7308 , \7310 );
mbuf \mul_7_15_g34273/U$1 ( \7312 , \5641 );
mnot \mul_7_15_g34184/U$3 ( \7313 , \7312 );
mbuf \mul_7_15_g34305/U$1 ( \7314 , \5706 );
mbuf \mul_7_15_g34283/U$1 ( \7315 , \5618 );
mand \mul_7_15_g34263/U$1 ( \7316 , \7314 , \7315 );
mnot \mul_7_15_g34192/U$3 ( \7317 , \7316 );
mnot \mul_7_15_g34198/U$2 ( \7318 , \7154 );
mnand \mul_7_15_g34210/U$1 ( \7319 , \6290 , \7137 );
mnand \mul_7_15_g34198/U$1 ( \7320 , \7318 , \7319 );
mnot \mul_7_15_g34192/U$4 ( \7321 , \7320 );
mor \mul_7_15_g34192/U$2 ( \7322 , \7317 , \7321 );
mbuf \mul_7_15_g34309/U$1 ( \7323 , \7159 );
mnot \mul_7_15_g34307/U$1 ( \7324 , \7323 );
mand \mul_7_15_g34248/U$2 ( \7325 , \7324 , \7315 );
mnot \mul_7_15_g34277/U$1 ( \7326 , \7160 );
mnor \mul_7_15_g34248/U$1 ( \7327 , \7325 , \7326 );
mnand \mul_7_15_g34192/U$1 ( \7328 , \7322 , \7327 );
mnot \mul_7_15_g34184/U$4 ( \7329 , \7328 );
mor \mul_7_15_g34184/U$2 ( \7330 , \7313 , \7329 );
mnand \mul_7_15_g34184/U$1 ( \7331 , \7330 , \7165 );
mnand \mul_7_15_g34243/U$1 ( \7332 , \7163 , \7167 );
mnot \mul_7_15_g34242/U$1 ( \7333 , \7332 );
mand \mul_7_15_g34180/U$2 ( \7334 , \7331 , \7333 );
mnot \mul_7_15_g34180/U$4 ( \7335 , \7331 );
mand \mul_7_15_g34180/U$3 ( \7336 , \7335 , \7332 );
mnor \mul_7_15_g34180/U$1 ( \7337 , \7334 , \7336 );
mnand \mul_7_15_g34311/U$1 ( \7338 , \7304 , \5004 );
mnot \mul_7_15_g34188/U$3 ( \7339 , \7338 );
mnot \mul_7_15_g34188/U$4 ( \7340 , \7241 );
mor \mul_7_15_g34188/U$2 ( \7341 , \7339 , \7340 );
mor \mul_7_15_g34188/U$5 ( \7342 , \7170 , \7338 );
mnand \mul_7_15_g34188/U$1 ( \7343 , \7341 , \7342 );
mnot \mul_7_15_g34193/U$3 ( \7344 , \7314 );
mbuf \fopt36714/U$1 ( \7345 , \7320 );
mnot \mul_7_15_g34193/U$4 ( \7346 , \7345 );
mor \mul_7_15_g34193/U$2 ( \7347 , \7344 , \7346 );
mnand \mul_7_15_g34193/U$1 ( \7348 , \7347 , \7323 );
mnand \mul_7_15_g34265/U$1 ( \7349 , \7160 , \7315 );
mnot \mul_7_15_g34264/U$1 ( \7350 , \7349 );
mand \mul_7_15_g34190/U$2 ( \7351 , \7348 , \7350 );
mnot \mul_7_15_g34190/U$4 ( \7352 , \7348 );
mand \mul_7_15_g34190/U$3 ( \7353 , \7352 , \7349 );
mnor \mul_7_15_g34190/U$1 ( \7354 , \7351 , \7353 );
mnand \mul_7_15_g34280/U$1 ( \7355 , \7323 , \7314 );
mnot \mul_7_15_g34279/U$1 ( \7356 , \7355 );
mand \mul_7_15_g34196/U$2 ( \7357 , \7345 , \7356 );
mnot \mul_7_15_g34196/U$4 ( \7358 , \7345 );
mand \mul_7_15_g34196/U$3 ( \7359 , \7358 , \7355 );
mnor \mul_7_15_g34196/U$1 ( \7360 , \7357 , \7359 );
mbuf \fopt36859/U$1 ( \7361 , \6034 );
mnot \mul_7_15_g34203/U$3 ( \7362 , \7361 );
mnot \mul_7_15_g34211/U$3 ( \7363 , \6279 );
mnot \mul_7_15_g34211/U$4 ( \7364 , \7137 );
mor \mul_7_15_g34211/U$2 ( \7365 , \7363 , \7364 );
mnand \mul_7_15_g34211/U$1 ( \7366 , \7365 , \7145 );
mnot \mul_7_15_g34203/U$4 ( \7367 , \7366 );
mor \mul_7_15_g34203/U$2 ( \7368 , \7362 , \7367 );
mnand \mul_7_15_g34203/U$1 ( \7369 , \7368 , \7147 );
mnand \mul_7_15_g34313/U$1 ( \7370 , \6288 , \7153 );
mnot \mul_7_15_g34312/U$1 ( \7371 , \7370 );
mand \mul_7_15_g34199/U$2 ( \7372 , \7369 , \7371 );
mnot \mul_7_15_g34199/U$4 ( \7373 , \7369 );
mand \mul_7_15_g34199/U$3 ( \7374 , \7373 , \7370 );
mnor \mul_7_15_g34199/U$1 ( \7375 , \7372 , \7374 );
mnand \mul_7_15_g34227/U$1 ( \7376 , \7147 , \7361 );
mnot \mul_7_15_g34226/U$1 ( \7377 , \7376 );
mand \mul_7_15_g34204/U$2 ( \7378 , \7366 , \7377 );
mnot \mul_7_15_g34204/U$4 ( \7379 , \7366 );
mand \mul_7_15_g34204/U$3 ( \7380 , \7379 , \7376 );
mnor \mul_7_15_g34204/U$1 ( \7381 , \7378 , \7380 );
mnot \mul_7_15_g34212/U$3 ( \7382 , \6278 );
mbuf \fopt36948/U$1 ( \7383 , \7137 );
mnot \mul_7_15_g34212/U$4 ( \7384 , \7383 );
mor \mul_7_15_g34212/U$2 ( \7385 , \7382 , \7384 );
mnand \mul_7_15_g34212/U$1 ( \7386 , \7385 , \7142 );
mnand \mul_7_15_g34229/U$1 ( \7387 , \6151 , \7140 );
mnot \mul_7_15_g34228/U$1 ( \7388 , \7387 );
mand \mul_7_15_g34205/U$2 ( \7389 , \7386 , \7388 );
mnot \mul_7_15_g34205/U$4 ( \7390 , \7386 );
mand \mul_7_15_g34205/U$3 ( \7391 , \7390 , \7387 );
mnor \mul_7_15_g34205/U$1 ( \7392 , \7389 , \7391 );
mnand \mul_7_15_g34245/U$1 ( \7393 , \7142 , \6278 );
mnot \mul_7_15_g34214/U$3 ( \7394 , \7393 );
mnot \mul_7_15_g34214/U$4 ( \7395 , \7383 );
mor \mul_7_15_g34214/U$2 ( \7396 , \7394 , \7395 );
mor \mul_7_15_g34214/U$5 ( \7397 , \7393 , \7383 );
mnand \mul_7_15_g34214/U$1 ( \7398 , \7396 , \7397 );
mbuf \mul_7_15_g34356/U$1 ( \7399 , \7068 );
mnot \mul_7_15_g34247/U$3 ( \7400 , \7399 );
mnot \mul_7_15_g34302/U$3 ( \7401 , \7115 );
mnot \mul_7_15_g34302/U$4 ( \7402 , \6983 );
mor \mul_7_15_g34302/U$2 ( \7403 , \7401 , \7402 );
mbuf \mul_7_15_fopt36299/U$1 ( \7404 , \7127 );
mnot \mul_7_15_g36437/U$2 ( \7405 , \7404 );
mnor \mul_7_15_g36437/U$1 ( \7406 , \7405 , \7124 );
mnand \mul_7_15_g34302/U$1 ( \7407 , \7403 , \7406 );
mnot \mul_7_15_g34247/U$4 ( \7408 , \7407 );
mor \mul_7_15_g34247/U$2 ( \7409 , \7400 , \7408 );
mnot \mul_7_15_g34361/U$1 ( \7410 , \7129 );
mnot \mul_7_15_g34360/U$1 ( \7411 , \7410 );
mnand \mul_7_15_g34247/U$1 ( \7412 , \7409 , \7411 );
mnand \mul_7_15_g34316/U$1 ( \7413 , \7119 , \7135 );
mnot \mul_7_15_g34315/U$1 ( \7414 , \7413 );
mand \mul_7_15_g34223/U$2 ( \7415 , \7412 , \7414 );
mnot \mul_7_15_g34223/U$4 ( \7416 , \7412 );
mand \mul_7_15_g34223/U$3 ( \7417 , \7416 , \7413 );
mnor \mul_7_15_g34223/U$1 ( \7418 , \7415 , \7417 );
mnand \mul_7_15_g34244/U$1 ( \7419 , \7165 , \7312 );
mnot \mul_7_15_g34327/U$2 ( \7420 , \7410 );
mnand \mul_7_15_g34327/U$1 ( \7421 , \7420 , \7399 );
mnot \mul_7_15_g34253/U$3 ( \7422 , \7421 );
mnot \mul_7_15_g34253/U$4 ( \7423 , \7407 );
mor \mul_7_15_g34253/U$2 ( \7424 , \7422 , \7423 );
mor \mul_7_15_g34253/U$5 ( \7425 , \7421 , \7407 );
mnand \mul_7_15_g34253/U$1 ( \7426 , \7424 , \7425 );
mnot \mul_7_15_g34286/U$3 ( \7427 , \7114 );
mnot \mul_7_15_g34286/U$4 ( \7428 , \6983 );
mor \mul_7_15_g34286/U$2 ( \7429 , \7427 , \7428 );
mnand \mul_7_15_g34286/U$1 ( \7430 , \7429 , \7123 );
mnand \mul_7_15_g34329/U$1 ( \7431 , \7404 , \7103 );
mnot \mul_7_15_g34328/U$1 ( \7432 , \7431 );
mand \mul_7_15_g34254/U$2 ( \7433 , \7430 , \7432 );
mnot \mul_7_15_g34254/U$4 ( \7434 , \7430 );
mand \mul_7_15_g34254/U$3 ( \7435 , \7434 , \7431 );
mnor \mul_7_15_g34254/U$1 ( \7436 , \7433 , \7435 );
mbuf \mul_7_15_g34458/U$1 ( \7437 , \6964 );
mnot \mul_7_15_g34287/U$3 ( \7438 , \7437 );
mnot \mul_7_15_g34347/U$3 ( \7439 , \6954 );
mnot \mul_7_15_g34347/U$4 ( \7440 , \6601 );
mor \mul_7_15_g34347/U$2 ( \7441 , \7439 , \7440 );
mnand \mul_7_15_g34460/U$1 ( \7442 , \6978 , \6944 );
mnand \mul_7_15_g34347/U$1 ( \7443 , \7441 , \7442 );
mnot \mul_7_15_g34287/U$4 ( \7444 , \7443 );
mor \mul_7_15_g34287/U$2 ( \7445 , \7438 , \7444 );
mnand \mul_7_15_g34287/U$1 ( \7446 , \7445 , \6973 );
mnand \mul_7_15_g34403/U$1 ( \7447 , \6981 , \6970 );
mnot \mul_7_15_g34402/U$1 ( \7448 , \7447 );
mand \mul_7_15_g34255/U$2 ( \7449 , \7446 , \7448 );
mnot \mul_7_15_g34255/U$4 ( \7450 , \7446 );
mand \mul_7_15_g34255/U$3 ( \7451 , \7450 , \7447 );
mnor \mul_7_15_g34255/U$1 ( \7452 , \7449 , \7451 );
mnand \mul_7_15_g34352/U$1 ( \7453 , \7114 , \7123 );
mnot \mul_7_15_g34293/U$3 ( \7454 , \7453 );
mnot \mul_7_15_g34293/U$4 ( \7455 , \6983 );
mor \mul_7_15_g34293/U$2 ( \7456 , \7454 , \7455 );
mor \mul_7_15_g34293/U$5 ( \7457 , \7453 , \6983 );
mnand \mul_7_15_g34293/U$1 ( \7458 , \7456 , \7457 );
mnand \mul_7_15_g34444/U$1 ( \7459 , \7437 , \6973 );
mnot \mul_7_15_g34443/U$1 ( \7460 , \7459 );
mand \mul_7_15_g34294/U$2 ( \7461 , \7443 , \7460 );
mnot \mul_7_15_g34294/U$4 ( \7462 , \7443 );
mand \mul_7_15_g34294/U$3 ( \7463 , \7462 , \7459 );
mnor \mul_7_15_g34294/U$1 ( \7464 , \7461 , \7463 );
mnot \mul_7_15_g34345/U$3 ( \7465 , \6953 );
mnot \mul_7_15_g34345/U$4 ( \7466 , \6601 );
mor \mul_7_15_g34345/U$2 ( \7467 , \7465 , \7466 );
mnand \mul_7_15_g34345/U$1 ( \7468 , \7467 , \6977 );
mnand \mul_7_15_g34486/U$1 ( \7469 , \6976 , \6944 );
mnot \mul_7_15_g34485/U$1 ( \7470 , \7469 );
mand \mul_7_15_g34295/U$2 ( \7471 , \7468 , \7470 );
mnot \mul_7_15_g34295/U$4 ( \7472 , \7468 );
mand \mul_7_15_g34295/U$3 ( \7473 , \7472 , \7469 );
mnor \mul_7_15_g34295/U$1 ( \7474 , \7471 , \7473 );
mnand \mul_7_15_g34523/U$1 ( \7475 , \6977 , \6953 );
mnot \mul_7_15_g34346/U$3 ( \7476 , \7475 );
mnot \mul_7_15_g34346/U$4 ( \7477 , \6601 );
mor \mul_7_15_g34346/U$2 ( \7478 , \7476 , \7477 );
mor \mul_7_15_g34346/U$5 ( \7479 , \7475 , \6601 );
mnand \mul_7_15_g34346/U$1 ( \7480 , \7478 , \7479 );
mxor \mul_7_15_g34389/U$1 ( \7481 , \6364 , \6428 );
mxor \mul_7_15_g34389/U$1_r1 ( \7482 , \7481 , \6598 );
mand \mul_7_15_g36379/U$1 ( \7483 , \6592 , \6589 );
mand \mul_7_15_g34536/U$2 ( \7484 , \7483 , \6571 );
mnot \mul_7_15_g34536/U$4 ( \7485 , \7483 );
mnot \mul_7_15_g34590/U$1 ( \7486 , \6571 );
mand \mul_7_15_g34536/U$3 ( \7487 , \7485 , \7486 );
mnor \mul_7_15_g34536/U$1 ( \7488 , \7484 , \7487 );
mnand \mul_7_15_g34575/U$1 ( \7489 , \6597 , \6471 );
mnot \mul_7_15_g34630/U$3 ( \7490 , \6567 );
mnand \mul_7_15_g34715/U$1 ( \7491 , \6570 , \6515 );
mnot \mul_7_15_g34630/U$4 ( \7492 , \7491 );
mor \mul_7_15_g34630/U$2 ( \7493 , \7490 , \7492 );
mor \mul_7_15_g34630/U$5 ( \7494 , \6567 , \7491 );
mnand \mul_7_15_g34630/U$1 ( \7495 , \7493 , \7494 );
mxor \mul_7_15_g34698/U$1 ( \7496 , \6526 , \6558 );
mxor \mul_7_15_g34698/U$1_r1 ( \7497 , \7496 , \6564 );
mnand \mul_7_15_g34995/U$1 ( \7498 , \6557 , \6539 );
mand \mul_7_15_g34885/U$2 ( \7499 , \7498 , \6552 );
mnot \mul_7_15_g34885/U$4 ( \7500 , \7498 );
mand \mul_7_15_g34885/U$3 ( \7501 , \7500 , \6553 );
mnor \mul_7_15_g34885/U$1 ( \7502 , \7499 , \7501 );
mnot \mul_7_15_g35007/U$2 ( \7503 , \6552 );
mnor \mul_7_15_g35009/U$1 ( \7504 , \6549 , \6551 );
mnor \mul_7_15_g35007/U$1 ( \7505 , \7503 , \7504 );
mnot \mul_7_15_g35784/U$1 ( \7506 , \6550 );
mxnor \mul_7_15_g36370/U$1 ( \7507 , \6593 , \7489 );
mxnor \g36456/U$1 ( \7508 , \7328 , \7419 );
endmodule

